module pure_cos_table(
     input              sclk,
     input              rst_n,
     output wire [15:0] pure_cos
    );
//
assign pure_cos[15:0] = cos_wave[15:0]; 
//
parameter lim = 999;
//
reg  [9:0] cnt;
reg [15:0] cos_wave;
//
always @(posedge sclk or negedge rst_n)
begin
     if (!rst_n)        cnt <= 0 ;
     else if (lim==cnt) cnt <= 0 ;
     else               cnt <= cnt+1 ; 
end
//
always @(posedge sclk or negedge rst_n)
begin
     if (!rst_n) cos_wave[15:0] = 16'h0000	;
     else
     case(cnt)
     0	: cos_wave[15:0] = 16'h7FFF	;
     1	: cos_wave[15:0] = 16'h7FFE	;
     2	: cos_wave[15:0] = 16'h7FFC	;
     3	: cos_wave[15:0] = 16'h7FF9	;
     4	: cos_wave[15:0] = 16'h7FF5	;
     5	: cos_wave[15:0] = 16'h7FEF	;
     6	: cos_wave[15:0] = 16'h7FE8	;
     7	: cos_wave[15:0] = 16'h7FDF	;
     8	: cos_wave[15:0] = 16'h7FD6	;
     9	: cos_wave[15:0] = 16'h7FCB	;
     10	: cos_wave[15:0] = 16'h7FBE	;
     11	: cos_wave[15:0] = 16'h7FB1	;
     12	: cos_wave[15:0] = 16'h7FA2	;
     13	: cos_wave[15:0] = 16'h7F92	;
     14	: cos_wave[15:0] = 16'h7F80	;
     15	: cos_wave[15:0] = 16'h7F6D	;
     16	: cos_wave[15:0] = 16'h7F59	;
     17	: cos_wave[15:0] = 16'h7F44	;
     18	: cos_wave[15:0] = 16'h7F2D	;
     19	: cos_wave[15:0] = 16'h7F15	;
     20	: cos_wave[15:0] = 16'h7EFC	;
     21	: cos_wave[15:0] = 16'h7EE2	;
     22	: cos_wave[15:0] = 16'h7EC6	;
     23	: cos_wave[15:0] = 16'h7EA9	;
     24	: cos_wave[15:0] = 16'h7E8A	;
     25	: cos_wave[15:0] = 16'h7E6B	;
     26	: cos_wave[15:0] = 16'h7E4A	;
     27	: cos_wave[15:0] = 16'h7E28	;
     28	: cos_wave[15:0] = 16'h7E04	;
     29	: cos_wave[15:0] = 16'h7DDF	;
     30	: cos_wave[15:0] = 16'h7DB9	;
     31	: cos_wave[15:0] = 16'h7D92	;
     32	: cos_wave[15:0] = 16'h7D6A	;
     33	: cos_wave[15:0] = 16'h7D40	;
     34	: cos_wave[15:0] = 16'h7D15	;
     35	: cos_wave[15:0] = 16'h7CE8	;
     36	: cos_wave[15:0] = 16'h7CBB	;
     37	: cos_wave[15:0] = 16'h7C8C	;
     38	: cos_wave[15:0] = 16'h7C5C	;
     39	: cos_wave[15:0] = 16'h7C2A	;
     40	: cos_wave[15:0] = 16'h7BF8	;
     41	: cos_wave[15:0] = 16'h7BC4	;
     42	: cos_wave[15:0] = 16'h7B8E	;
     43	: cos_wave[15:0] = 16'h7B58	;
     44	: cos_wave[15:0] = 16'h7B20	;
     45	: cos_wave[15:0] = 16'h7AE7	;
     46	: cos_wave[15:0] = 16'h7AAD	;
     47	: cos_wave[15:0] = 16'h7A72	;
     48	: cos_wave[15:0] = 16'h7A35	;
     49	: cos_wave[15:0] = 16'h79F7	;
     50	: cos_wave[15:0] = 16'h79B8	;
     51	: cos_wave[15:0] = 16'h7978	;
     52	: cos_wave[15:0] = 16'h7936	;
     53	: cos_wave[15:0] = 16'h78F3	;
     54	: cos_wave[15:0] = 16'h78AF	;
     55	: cos_wave[15:0] = 16'h786A	;
     56	: cos_wave[15:0] = 16'h7824	;
     57	: cos_wave[15:0] = 16'h77DC	;
     58	: cos_wave[15:0] = 16'h7793	;
     59	: cos_wave[15:0] = 16'h7749	;
     60	: cos_wave[15:0] = 16'h76FD	;
     61	: cos_wave[15:0] = 16'h76B1	;
     62	: cos_wave[15:0] = 16'h7663	;
     63	: cos_wave[15:0] = 16'h7614	;
     64	: cos_wave[15:0] = 16'h75C4	;
     65	: cos_wave[15:0] = 16'h7573	;
     66	: cos_wave[15:0] = 16'h7520	;
     67	: cos_wave[15:0] = 16'h74CD	;
     68	: cos_wave[15:0] = 16'h7478	;
     69	: cos_wave[15:0] = 16'h7422	;
     70	: cos_wave[15:0] = 16'h73CA	;
     71	: cos_wave[15:0] = 16'h7372	;
     72	: cos_wave[15:0] = 16'h7318	;
     73	: cos_wave[15:0] = 16'h72BE	;
     74	: cos_wave[15:0] = 16'h7262	;
     75	: cos_wave[15:0] = 16'h7205	;
     76	: cos_wave[15:0] = 16'h71A6	;
     77	: cos_wave[15:0] = 16'h7147	;
     78	: cos_wave[15:0] = 16'h70E6	;
     79	: cos_wave[15:0] = 16'h7085	;
     80	: cos_wave[15:0] = 16'h7022	;
     81	: cos_wave[15:0] = 16'h6FBE	;
     82	: cos_wave[15:0] = 16'h6F59	;
     83	: cos_wave[15:0] = 16'h6EF3	;
     84	: cos_wave[15:0] = 16'h6E8B	;
     85	: cos_wave[15:0] = 16'h6E23	;
     86	: cos_wave[15:0] = 16'h6DB9	;
     87	: cos_wave[15:0] = 16'h6D4F	;
     88	: cos_wave[15:0] = 16'h6CE3	;
     89	: cos_wave[15:0] = 16'h6C76	;
     90	: cos_wave[15:0] = 16'h6C08	;
     91	: cos_wave[15:0] = 16'h6B99	;
     92	: cos_wave[15:0] = 16'h6B29	;
     93	: cos_wave[15:0] = 16'h6AB8	;
     94	: cos_wave[15:0] = 16'h6A45	;
     95	: cos_wave[15:0] = 16'h69D2	;
     96	: cos_wave[15:0] = 16'h695D	;
     97	: cos_wave[15:0] = 16'h68E8	;
     98	: cos_wave[15:0] = 16'h6871	;
     99	: cos_wave[15:0] = 16'h67FA	;
     100: cos_wave[15:0] = 16'h6781	;
     101: cos_wave[15:0] = 16'h6707	;
     102: cos_wave[15:0] = 16'h668C	;
     103: cos_wave[15:0] = 16'h6611	;
     104: cos_wave[15:0] = 16'h6594	;
     105: cos_wave[15:0] = 16'h6516	;
     106: cos_wave[15:0] = 16'h6497	;
     107: cos_wave[15:0] = 16'h6417	;
     108: cos_wave[15:0] = 16'h6396	;
     109: cos_wave[15:0] = 16'h6314	;
     110: cos_wave[15:0] = 16'h6291	;
     111: cos_wave[15:0] = 16'h620D	;
     112: cos_wave[15:0] = 16'h6188	;
     113: cos_wave[15:0] = 16'h6102	;
     114: cos_wave[15:0] = 16'h607B	;
     115: cos_wave[15:0] = 16'h5FF3	;
     116: cos_wave[15:0] = 16'h5F6A	;
     117: cos_wave[15:0] = 16'h5EE0	;
     118: cos_wave[15:0] = 16'h5E56	;
     119: cos_wave[15:0] = 16'h5DCA	;
     120: cos_wave[15:0] = 16'h5D3D	;
     121: cos_wave[15:0] = 16'h5CB0	;
     122: cos_wave[15:0] = 16'h5C21	;
     123: cos_wave[15:0] = 16'h5B91	;
     124: cos_wave[15:0] = 16'h5B01	;
     125: cos_wave[15:0] = 16'h5A70	;
     126: cos_wave[15:0] = 16'h59DD	;
     127: cos_wave[15:0] = 16'h594A	;
     128: cos_wave[15:0] = 16'h58B6	;
     129: cos_wave[15:0] = 16'h5821	;
     130: cos_wave[15:0] = 16'h578B	;
     131: cos_wave[15:0] = 16'h56F4	;
     132: cos_wave[15:0] = 16'h565D	;
     133: cos_wave[15:0] = 16'h55C4	;
     134: cos_wave[15:0] = 16'h552B	;
     135: cos_wave[15:0] = 16'h5490	;
     136: cos_wave[15:0] = 16'h53F5	;
     137: cos_wave[15:0] = 16'h5359	;
     138: cos_wave[15:0] = 16'h52BC	;
     139: cos_wave[15:0] = 16'h521F	;
     140: cos_wave[15:0] = 16'h5180	;
     141: cos_wave[15:0] = 16'h50E1	;
     142: cos_wave[15:0] = 16'h5041	;
     143: cos_wave[15:0] = 16'h4FA0	;
     144: cos_wave[15:0] = 16'h4EFE	;
     145: cos_wave[15:0] = 16'h4E5C	;
     146: cos_wave[15:0] = 16'h4DB8	;
     147: cos_wave[15:0] = 16'h4D14	;
     148: cos_wave[15:0] = 16'h4C6F	;
     149: cos_wave[15:0] = 16'h4BC9	;
     150: cos_wave[15:0] = 16'h4B23	;
     151: cos_wave[15:0] = 16'h4A7C	;
     152: cos_wave[15:0] = 16'h49D4	;
     153: cos_wave[15:0] = 16'h492B	;
     154: cos_wave[15:0] = 16'h4882	;
     155: cos_wave[15:0] = 16'h47D7	;
     156: cos_wave[15:0] = 16'h472C	;
     157: cos_wave[15:0] = 16'h4681	;
     158: cos_wave[15:0] = 16'h45D4	;
     159: cos_wave[15:0] = 16'h4527	;
     160: cos_wave[15:0] = 16'h447A	;
     161: cos_wave[15:0] = 16'h43CB	;
     162: cos_wave[15:0] = 16'h431C	;
     163: cos_wave[15:0] = 16'h426C	;
     164: cos_wave[15:0] = 16'h41BC	;
     165: cos_wave[15:0] = 16'h410A	;
     166: cos_wave[15:0] = 16'h4059	;
     167: cos_wave[15:0] = 16'h3FA6	;
     168: cos_wave[15:0] = 16'h3EF3	;
     169: cos_wave[15:0] = 16'h3E3F	;
     170: cos_wave[15:0] = 16'h3D8B	;
     171: cos_wave[15:0] = 16'h3CD6	;
     172: cos_wave[15:0] = 16'h3C20	;
     173: cos_wave[15:0] = 16'h3B6A	;
     174: cos_wave[15:0] = 16'h3AB3	;
     175: cos_wave[15:0] = 16'h39FC	;
     176: cos_wave[15:0] = 16'h3944	;
     177: cos_wave[15:0] = 16'h388B	;
     178: cos_wave[15:0] = 16'h37D2	;
     179: cos_wave[15:0] = 16'h3718	;
     180: cos_wave[15:0] = 16'h365E	;
     181: cos_wave[15:0] = 16'h35A3	;
     182: cos_wave[15:0] = 16'h34E8	;
     183: cos_wave[15:0] = 16'h342C	;
     184: cos_wave[15:0] = 16'h336F	;
     185: cos_wave[15:0] = 16'h32B2	;
     186: cos_wave[15:0] = 16'h31F5	;
     187: cos_wave[15:0] = 16'h3137	;
     188: cos_wave[15:0] = 16'h3078	;
     189: cos_wave[15:0] = 16'h2FB9	;
     190: cos_wave[15:0] = 16'h2EFA	;
     191: cos_wave[15:0] = 16'h2E3A	;
     192: cos_wave[15:0] = 16'h2D7A	;
     193: cos_wave[15:0] = 16'h2CB9	;
     194: cos_wave[15:0] = 16'h2BF7	;
     195: cos_wave[15:0] = 16'h2B36	;
     196: cos_wave[15:0] = 16'h2A73	;
     197: cos_wave[15:0] = 16'h29B1	;
     198: cos_wave[15:0] = 16'h28EE	;
     199: cos_wave[15:0] = 16'h282A	;
     200: cos_wave[15:0] = 16'h2766	;
     201: cos_wave[15:0] = 16'h26A2	;
     202: cos_wave[15:0] = 16'h25DD	;
     203: cos_wave[15:0] = 16'h2518	;
     204: cos_wave[15:0] = 16'h2453	;
     205: cos_wave[15:0] = 16'h238D	;
     206: cos_wave[15:0] = 16'h22C7	;
     207: cos_wave[15:0] = 16'h2200	;
     208: cos_wave[15:0] = 16'h213A	;
     209: cos_wave[15:0] = 16'h2072	;
     210: cos_wave[15:0] = 16'h1FAB	;
     211: cos_wave[15:0] = 16'h1EE3	;
     212: cos_wave[15:0] = 16'h1E1B	;
     213: cos_wave[15:0] = 16'h1D52	;
     214: cos_wave[15:0] = 16'h1C8A	;
     215: cos_wave[15:0] = 16'h1BC1	;
     216: cos_wave[15:0] = 16'h1AF7	;
     217: cos_wave[15:0] = 16'h1A2E	;
     218: cos_wave[15:0] = 16'h1964	;
     219: cos_wave[15:0] = 16'h189A	;
     220: cos_wave[15:0] = 16'h17CF	;
     221: cos_wave[15:0] = 16'h1705	;
     222: cos_wave[15:0] = 16'h163A	;
     223: cos_wave[15:0] = 16'h156F	;
     224: cos_wave[15:0] = 16'h14A4	;
     225: cos_wave[15:0] = 16'h13D8	;
     226: cos_wave[15:0] = 16'h130C	;
     227: cos_wave[15:0] = 16'h1241	;
     228: cos_wave[15:0] = 16'h1174	;
     229: cos_wave[15:0] = 16'h10A8	;
     230: cos_wave[15:0] = 16'h0FDC	;
     231: cos_wave[15:0] = 16'h0F0F	;
     232: cos_wave[15:0] = 16'h0E42	;
     233: cos_wave[15:0] = 16'h0D76	;
     234: cos_wave[15:0] = 16'h0CA9	;
     235: cos_wave[15:0] = 16'h0BDB	;
     236: cos_wave[15:0] = 16'h0B0E	;
     237: cos_wave[15:0] = 16'h0A41	;
     238: cos_wave[15:0] = 16'h0973	;
     239: cos_wave[15:0] = 16'h08A6	;
     240: cos_wave[15:0] = 16'h07D8	;
     241: cos_wave[15:0] = 16'h070A	;
     242: cos_wave[15:0] = 16'h063D	;
     243: cos_wave[15:0] = 16'h056F	;
     244: cos_wave[15:0] = 16'h04A1	;
     245: cos_wave[15:0] = 16'h03D3	;
     246: cos_wave[15:0] = 16'h0305	;
     247: cos_wave[15:0] = 16'h0237	;
     248: cos_wave[15:0] = 16'h0169	;
     249: cos_wave[15:0] = 16'h009B	;
     250: cos_wave[15:0] = 16'hFFCC	;
     251: cos_wave[15:0] = 16'hFEFE	;
     252: cos_wave[15:0] = 16'hFE30	;
     253: cos_wave[15:0] = 16'hFD62	;
     254: cos_wave[15:0] = 16'hFC94	;
     255: cos_wave[15:0] = 16'hFBC6	;
     256: cos_wave[15:0] = 16'hFAF8	;
     257: cos_wave[15:0] = 16'hFA2A	;
     258: cos_wave[15:0] = 16'hF95D	;
     259: cos_wave[15:0] = 16'hF88F	;
     260: cos_wave[15:0] = 16'hF7C1	;
     261: cos_wave[15:0] = 16'hF6F3	;
     262: cos_wave[15:0] = 16'hF626	;
     263: cos_wave[15:0] = 16'hF559	;
     264: cos_wave[15:0] = 16'hF48B	;
     265: cos_wave[15:0] = 16'hF3BE	;
     266: cos_wave[15:0] = 16'hF2F1	;
     267: cos_wave[15:0] = 16'hF224	;
     268: cos_wave[15:0] = 16'hF157	;
     269: cos_wave[15:0] = 16'hF08B	;
     270: cos_wave[15:0] = 16'hEFBE	;
     271: cos_wave[15:0] = 16'hEEF2	;
     272: cos_wave[15:0] = 16'hEE26	;
     273: cos_wave[15:0] = 16'hED5A	;
     274: cos_wave[15:0] = 16'hEC8E	;
     275: cos_wave[15:0] = 16'hEBC2	;
     276: cos_wave[15:0] = 16'hEAF7	;
     277: cos_wave[15:0] = 16'hEA2C	;
     278: cos_wave[15:0] = 16'hE961	;
     279: cos_wave[15:0] = 16'hE896	;
     280: cos_wave[15:0] = 16'hE7CB	;
     281: cos_wave[15:0] = 16'hE701	;
     282: cos_wave[15:0] = 16'hE637	;
     283: cos_wave[15:0] = 16'hE56D	;
     284: cos_wave[15:0] = 16'hE4A4	;
     285: cos_wave[15:0] = 16'hE3DB	;
     286: cos_wave[15:0] = 16'hE312	;
     287: cos_wave[15:0] = 16'hE249	;
     288: cos_wave[15:0] = 16'hE181	;
     289: cos_wave[15:0] = 16'hE0B9	;
     290: cos_wave[15:0] = 16'hDFF1	;
     291: cos_wave[15:0] = 16'hDF2A	;
     292: cos_wave[15:0] = 16'hDE63	;
     293: cos_wave[15:0] = 16'hDD9C	;
     294: cos_wave[15:0] = 16'hDCD6	;
     295: cos_wave[15:0] = 16'hDC10	;
     296: cos_wave[15:0] = 16'hDB4A	;
     297: cos_wave[15:0] = 16'hDA85	;
     298: cos_wave[15:0] = 16'hD9C0	;
     299: cos_wave[15:0] = 16'hD8FC	;
     300: cos_wave[15:0] = 16'hD838	;
     301: cos_wave[15:0] = 16'hD774	;
     302: cos_wave[15:0] = 16'hD6B1	;
     303: cos_wave[15:0] = 16'hD5EE	;
     304: cos_wave[15:0] = 16'hD52B	;
     305: cos_wave[15:0] = 16'hD469	;
     306: cos_wave[15:0] = 16'hD3A8	;
     307: cos_wave[15:0] = 16'hD2E7	;
     308: cos_wave[15:0] = 16'hD226	;
     309: cos_wave[15:0] = 16'hD166	;
     310: cos_wave[15:0] = 16'hD0A6	;
     311: cos_wave[15:0] = 16'hCFE7	;
     312: cos_wave[15:0] = 16'hCF28	;
     313: cos_wave[15:0] = 16'hCE6A	;
     314: cos_wave[15:0] = 16'hCDAC	;
     315: cos_wave[15:0] = 16'hCCEF	;
     316: cos_wave[15:0] = 16'hCC32	;
     317: cos_wave[15:0] = 16'hCB76	;
     318: cos_wave[15:0] = 16'hCABB	;
     319: cos_wave[15:0] = 16'hC9FF	;
     320: cos_wave[15:0] = 16'hC945	;
     321: cos_wave[15:0] = 16'hC88B	;
     322: cos_wave[15:0] = 16'hC7D1	;
     323: cos_wave[15:0] = 16'hC718	;
     324: cos_wave[15:0] = 16'hC660	;
     325: cos_wave[15:0] = 16'hC5A8	;
     326: cos_wave[15:0] = 16'hC4F1	;
     327: cos_wave[15:0] = 16'hC43B	;
     328: cos_wave[15:0] = 16'hC385	;
     329: cos_wave[15:0] = 16'hC2D0	;
     330: cos_wave[15:0] = 16'hC21B	;
     331: cos_wave[15:0] = 16'hC167	;
     332: cos_wave[15:0] = 16'hC0B3	;
     333: cos_wave[15:0] = 16'hC000	;
     334: cos_wave[15:0] = 16'hBF4E	;
     335: cos_wave[15:0] = 16'hBE9D	;
     336: cos_wave[15:0] = 16'hBDEC	;
     337: cos_wave[15:0] = 16'hBD3C	;
     338: cos_wave[15:0] = 16'hBC8C	;
     339: cos_wave[15:0] = 16'hBBDE	;
     340: cos_wave[15:0] = 16'hBB2F	;
     341: cos_wave[15:0] = 16'hBA82	;
     342: cos_wave[15:0] = 16'hB9D5	;
     343: cos_wave[15:0] = 16'hB929	;
     344: cos_wave[15:0] = 16'hB87E	;
     345: cos_wave[15:0] = 16'hB7D3	;
     346: cos_wave[15:0] = 16'hB72A	;
     347: cos_wave[15:0] = 16'hB681	;
     348: cos_wave[15:0] = 16'hB5D8	;
     349: cos_wave[15:0] = 16'hB531	;
     350: cos_wave[15:0] = 16'hB48A	;
     351: cos_wave[15:0] = 16'hB3E4	;
     352: cos_wave[15:0] = 16'hB33E	;
     353: cos_wave[15:0] = 16'hB29A	;
     354: cos_wave[15:0] = 16'hB1F6	;
     355: cos_wave[15:0] = 16'hB153	;
     356: cos_wave[15:0] = 16'hB0B1	;
     357: cos_wave[15:0] = 16'hB010	;
     358: cos_wave[15:0] = 16'hAF6F	;
     359: cos_wave[15:0] = 16'hAECF	;
     360: cos_wave[15:0] = 16'hAE30	;
     361: cos_wave[15:0] = 16'hAD92	;
     362: cos_wave[15:0] = 16'hACF5	;
     363: cos_wave[15:0] = 16'hAC59	;
     364: cos_wave[15:0] = 16'hABBD	;
     365: cos_wave[15:0] = 16'hAB22	;
     366: cos_wave[15:0] = 16'hAA89	;
     367: cos_wave[15:0] = 16'hA9F0	;
     368: cos_wave[15:0] = 16'hA957	;
     369: cos_wave[15:0] = 16'hA8C0	;
     370: cos_wave[15:0] = 16'hA82A	;
     371: cos_wave[15:0] = 16'hA794	;
     372: cos_wave[15:0] = 16'hA700	;
     373: cos_wave[15:0] = 16'hA66C	;
     374: cos_wave[15:0] = 16'hA5D9	;
     375: cos_wave[15:0] = 16'hA548	;
     376: cos_wave[15:0] = 16'hA4B7	;
     377: cos_wave[15:0] = 16'hA427	;
     378: cos_wave[15:0] = 16'hA398	;
     379: cos_wave[15:0] = 16'hA30A	;
     380: cos_wave[15:0] = 16'hA27C	;
     381: cos_wave[15:0] = 16'hA1F0	;
     382: cos_wave[15:0] = 16'hA165	;
     383: cos_wave[15:0] = 16'hA0DA	;
     384: cos_wave[15:0] = 16'hA051	;
     385: cos_wave[15:0] = 16'h9FC9	;
     386: cos_wave[15:0] = 16'h9F41	;
     387: cos_wave[15:0] = 16'h9EBB	;
     388: cos_wave[15:0] = 16'h9E35	;
     389: cos_wave[15:0] = 16'h9DB1	;
     390: cos_wave[15:0] = 16'h9D2D	;
     391: cos_wave[15:0] = 16'h9CAB	;
     392: cos_wave[15:0] = 16'h9C29	;
     393: cos_wave[15:0] = 16'h9BA9	;
     394: cos_wave[15:0] = 16'h9B2A	;
     395: cos_wave[15:0] = 16'h9AAB	;
     396: cos_wave[15:0] = 16'h9A2E	;
     397: cos_wave[15:0] = 16'h99B1	;
     398: cos_wave[15:0] = 16'h9936	;
     399: cos_wave[15:0] = 16'h98BC	;
     400: cos_wave[15:0] = 16'h9843	;
     401: cos_wave[15:0] = 16'h97CA	;
     402: cos_wave[15:0] = 16'h9753	;
     403: cos_wave[15:0] = 16'h96DD	;
     404: cos_wave[15:0] = 16'h9668	;
     405: cos_wave[15:0] = 16'h95F4	;
     406: cos_wave[15:0] = 16'h9581	;
     407: cos_wave[15:0] = 16'h9510	;
     408: cos_wave[15:0] = 16'h949F	;
     409: cos_wave[15:0] = 16'h942F	;
     410: cos_wave[15:0] = 16'h93C1	;
     411: cos_wave[15:0] = 16'h9353	;
     412: cos_wave[15:0] = 16'h92E7	;
     413: cos_wave[15:0] = 16'h927C	;
     414: cos_wave[15:0] = 16'h9212	;
     415: cos_wave[15:0] = 16'h91A9	;
     416: cos_wave[15:0] = 16'h9141	;
     417: cos_wave[15:0] = 16'h90DA	;
     418: cos_wave[15:0] = 16'h9074	;
     419: cos_wave[15:0] = 16'h9010	;
     420: cos_wave[15:0] = 16'h8FAC	;
     421: cos_wave[15:0] = 16'h8F4A	;
     422: cos_wave[15:0] = 16'h8EE9	;
     423: cos_wave[15:0] = 16'h8E89	;
     424: cos_wave[15:0] = 16'h8E2A	;
     425: cos_wave[15:0] = 16'h8DCD	;
     426: cos_wave[15:0] = 16'h8D70	;
     427: cos_wave[15:0] = 16'h8D15	;
     428: cos_wave[15:0] = 16'h8CBB	;
     429: cos_wave[15:0] = 16'h8C62	;
     430: cos_wave[15:0] = 16'h8C0A	;
     431: cos_wave[15:0] = 16'h8BB3	;
     432: cos_wave[15:0] = 16'h8B5E	;
     433: cos_wave[15:0] = 16'h8B09	;
     434: cos_wave[15:0] = 16'h8AB6	;
     435: cos_wave[15:0] = 16'h8A64	;
     436: cos_wave[15:0] = 16'h8A14	;
     437: cos_wave[15:0] = 16'h89C4	;
     438: cos_wave[15:0] = 16'h8976	;
     439: cos_wave[15:0] = 16'h8929	;
     440: cos_wave[15:0] = 16'h88DD	;
     441: cos_wave[15:0] = 16'h8892	;
     442: cos_wave[15:0] = 16'h8848	;
     443: cos_wave[15:0] = 16'h8800	;
     444: cos_wave[15:0] = 16'h87B9	;
     445: cos_wave[15:0] = 16'h8773	;
     446: cos_wave[15:0] = 16'h872F	;
     447: cos_wave[15:0] = 16'h86EB	;
     448: cos_wave[15:0] = 16'h86A9	;
     449: cos_wave[15:0] = 16'h8668	;
     450: cos_wave[15:0] = 16'h8628	;
     451: cos_wave[15:0] = 16'h85EA	;
     452: cos_wave[15:0] = 16'h85AC	;
     453: cos_wave[15:0] = 16'h8570	;
     454: cos_wave[15:0] = 16'h8536	;
     455: cos_wave[15:0] = 16'h84FC	;
     456: cos_wave[15:0] = 16'h84C4	;
     457: cos_wave[15:0] = 16'h848D	;
     458: cos_wave[15:0] = 16'h8457	;
     459: cos_wave[15:0] = 16'h8422	;
     460: cos_wave[15:0] = 16'h83EF	;
     461: cos_wave[15:0] = 16'h83BD	;
     462: cos_wave[15:0] = 16'h838C	;
     463: cos_wave[15:0] = 16'h835D	;
     464: cos_wave[15:0] = 16'h832E	;
     465: cos_wave[15:0] = 16'h8301	;
     466: cos_wave[15:0] = 16'h82D6	;
     467: cos_wave[15:0] = 16'h82AB	;
     468: cos_wave[15:0] = 16'h8282	;
     469: cos_wave[15:0] = 16'h825A	;
     470: cos_wave[15:0] = 16'h8233	;
     471: cos_wave[15:0] = 16'h820E	;
     472: cos_wave[15:0] = 16'h81EA	;
     473: cos_wave[15:0] = 16'h81C7	;
     474: cos_wave[15:0] = 16'h81A6	;
     475: cos_wave[15:0] = 16'h8185	;
     476: cos_wave[15:0] = 16'h8166	;
     477: cos_wave[15:0] = 16'h8149	;
     478: cos_wave[15:0] = 16'h812C	;
     479: cos_wave[15:0] = 16'h8111	;
     480: cos_wave[15:0] = 16'h80F7	;
     481: cos_wave[15:0] = 16'h80DF	;
     482: cos_wave[15:0] = 16'h80C7	;
     483: cos_wave[15:0] = 16'h80B1	;
     484: cos_wave[15:0] = 16'h809D	;
     485: cos_wave[15:0] = 16'h8089	;
     486: cos_wave[15:0] = 16'h8077	;
     487: cos_wave[15:0] = 16'h8066	;
     488: cos_wave[15:0] = 16'h8057	;
     489: cos_wave[15:0] = 16'h8048	;
     490: cos_wave[15:0] = 16'h803B	;
     491: cos_wave[15:0] = 16'h8030	;
     492: cos_wave[15:0] = 16'h8025	;
     493: cos_wave[15:0] = 16'h801C	;
     494: cos_wave[15:0] = 16'h8015	;
     495: cos_wave[15:0] = 16'h800E	;
     496: cos_wave[15:0] = 16'h8009	;
     497: cos_wave[15:0] = 16'h8005	;
     498: cos_wave[15:0] = 16'h8002	;
     499: cos_wave[15:0] = 16'h8001	;
     500: cos_wave[15:0] = 16'h8001	;
     501: cos_wave[15:0] = 16'h8002	;
     502: cos_wave[15:0] = 16'h8005	;
     503: cos_wave[15:0] = 16'h8009	;
     504: cos_wave[15:0] = 16'h800E	;
     505: cos_wave[15:0] = 16'h8015	;
     506: cos_wave[15:0] = 16'h801C	;
     507: cos_wave[15:0] = 16'h8025	;
     508: cos_wave[15:0] = 16'h8030	;
     509: cos_wave[15:0] = 16'h803B	;
     510: cos_wave[15:0] = 16'h8048	;
     511: cos_wave[15:0] = 16'h8057	;
     512: cos_wave[15:0] = 16'h8066	;
     513: cos_wave[15:0] = 16'h8077	;
     514: cos_wave[15:0] = 16'h8089	;
     515: cos_wave[15:0] = 16'h809D	;
     516: cos_wave[15:0] = 16'h80B1	;
     517: cos_wave[15:0] = 16'h80C7	;
     518: cos_wave[15:0] = 16'h80DF	;
     519: cos_wave[15:0] = 16'h80F7	;
     520: cos_wave[15:0] = 16'h8111	;
     521: cos_wave[15:0] = 16'h812C	;
     522: cos_wave[15:0] = 16'h8149	;
     523: cos_wave[15:0] = 16'h8166	;
     524: cos_wave[15:0] = 16'h8185	;
     525: cos_wave[15:0] = 16'h81A6	;
     526: cos_wave[15:0] = 16'h81C7	;
     527: cos_wave[15:0] = 16'h81EA	;
     528: cos_wave[15:0] = 16'h820E	;
     529: cos_wave[15:0] = 16'h8233	;
     530: cos_wave[15:0] = 16'h825A	;
     531: cos_wave[15:0] = 16'h8282	;
     532: cos_wave[15:0] = 16'h82AB	;
     533: cos_wave[15:0] = 16'h82D6	;
     534: cos_wave[15:0] = 16'h8301	;
     535: cos_wave[15:0] = 16'h832E	;
     536: cos_wave[15:0] = 16'h835D	;
     537: cos_wave[15:0] = 16'h838C	;
     538: cos_wave[15:0] = 16'h83BD	;
     539: cos_wave[15:0] = 16'h83EF	;
     540: cos_wave[15:0] = 16'h8422	;
     541: cos_wave[15:0] = 16'h8457	;
     542: cos_wave[15:0] = 16'h848D	;
     543: cos_wave[15:0] = 16'h84C4	;
     544: cos_wave[15:0] = 16'h84FC	;
     545: cos_wave[15:0] = 16'h8536	;
     546: cos_wave[15:0] = 16'h8570	;
     547: cos_wave[15:0] = 16'h85AC	;
     548: cos_wave[15:0] = 16'h85EA	;
     549: cos_wave[15:0] = 16'h8628	;
     550: cos_wave[15:0] = 16'h8668	;
     551: cos_wave[15:0] = 16'h86A9	;
     552: cos_wave[15:0] = 16'h86EB	;
     553: cos_wave[15:0] = 16'h872F	;
     554: cos_wave[15:0] = 16'h8773	;
     555: cos_wave[15:0] = 16'h87B9	;
     556: cos_wave[15:0] = 16'h8800	;
     557: cos_wave[15:0] = 16'h8848	;
     558: cos_wave[15:0] = 16'h8892	;
     559: cos_wave[15:0] = 16'h88DD	;
     560: cos_wave[15:0] = 16'h8929	;
     561: cos_wave[15:0] = 16'h8976	;
     562: cos_wave[15:0] = 16'h89C4	;
     563: cos_wave[15:0] = 16'h8A14	;
     564: cos_wave[15:0] = 16'h8A64	;
     565: cos_wave[15:0] = 16'h8AB6	;
     566: cos_wave[15:0] = 16'h8B09	;
     567: cos_wave[15:0] = 16'h8B5E	;
     568: cos_wave[15:0] = 16'h8BB3	;
     569: cos_wave[15:0] = 16'h8C0A	;
     570: cos_wave[15:0] = 16'h8C62	;
     571: cos_wave[15:0] = 16'h8CBB	;
     572: cos_wave[15:0] = 16'h8D15	;
     573: cos_wave[15:0] = 16'h8D70	;
     574: cos_wave[15:0] = 16'h8DCD	;
     575: cos_wave[15:0] = 16'h8E2A	;
     576: cos_wave[15:0] = 16'h8E89	;
     577: cos_wave[15:0] = 16'h8EE9	;
     578: cos_wave[15:0] = 16'h8F4A	;
     579: cos_wave[15:0] = 16'h8FAC	;
     580: cos_wave[15:0] = 16'h9010	;
     581: cos_wave[15:0] = 16'h9074	;
     582: cos_wave[15:0] = 16'h90DA	;
     583: cos_wave[15:0] = 16'h9141	;
     584: cos_wave[15:0] = 16'h91A9	;
     585: cos_wave[15:0] = 16'h9212	;
     586: cos_wave[15:0] = 16'h927C	;
     587: cos_wave[15:0] = 16'h92E7	;
     588: cos_wave[15:0] = 16'h9353	;
     589: cos_wave[15:0] = 16'h93C1	;
     590: cos_wave[15:0] = 16'h942F	;
     591: cos_wave[15:0] = 16'h949F	;
     592: cos_wave[15:0] = 16'h9510	;
     593: cos_wave[15:0] = 16'h9581	;
     594: cos_wave[15:0] = 16'h95F4	;
     595: cos_wave[15:0] = 16'h9668	;
     596: cos_wave[15:0] = 16'h96DD	;
     597: cos_wave[15:0] = 16'h9753	;
     598: cos_wave[15:0] = 16'h97CA	;
     599: cos_wave[15:0] = 16'h9843	;
     600: cos_wave[15:0] = 16'h98BC	;
     601: cos_wave[15:0] = 16'h9936	;
     602: cos_wave[15:0] = 16'h99B1	;
     603: cos_wave[15:0] = 16'h9A2E	;
     604: cos_wave[15:0] = 16'h9AAB	;
     605: cos_wave[15:0] = 16'h9B2A	;
     606: cos_wave[15:0] = 16'h9BA9	;
     607: cos_wave[15:0] = 16'h9C29	;
     608: cos_wave[15:0] = 16'h9CAB	;
     609: cos_wave[15:0] = 16'h9D2D	;
     610: cos_wave[15:0] = 16'h9DB1	;
     611: cos_wave[15:0] = 16'h9E35	;
     612: cos_wave[15:0] = 16'h9EBB	;
     613: cos_wave[15:0] = 16'h9F41	;
     614: cos_wave[15:0] = 16'h9FC9	;
     615: cos_wave[15:0] = 16'hA051	;
     616: cos_wave[15:0] = 16'hA0DA	;
     617: cos_wave[15:0] = 16'hA165	;
     618: cos_wave[15:0] = 16'hA1F0	;
     619: cos_wave[15:0] = 16'hA27C	;
     620: cos_wave[15:0] = 16'hA30A	;
     621: cos_wave[15:0] = 16'hA398	;
     622: cos_wave[15:0] = 16'hA427	;
     623: cos_wave[15:0] = 16'hA4B7	;
     624: cos_wave[15:0] = 16'hA548	;
     625: cos_wave[15:0] = 16'hA5D9	;
     626: cos_wave[15:0] = 16'hA66C	;
     627: cos_wave[15:0] = 16'hA700	;
     628: cos_wave[15:0] = 16'hA794	;
     629: cos_wave[15:0] = 16'hA82A	;
     630: cos_wave[15:0] = 16'hA8C0	;
     631: cos_wave[15:0] = 16'hA957	;
     632: cos_wave[15:0] = 16'hA9F0	;
     633: cos_wave[15:0] = 16'hAA89	;
     634: cos_wave[15:0] = 16'hAB22	;
     635: cos_wave[15:0] = 16'hABBD	;
     636: cos_wave[15:0] = 16'hAC59	;
     637: cos_wave[15:0] = 16'hACF5	;
     638: cos_wave[15:0] = 16'hAD92	;
     639: cos_wave[15:0] = 16'hAE30	;
     640: cos_wave[15:0] = 16'hAECF	;
     641: cos_wave[15:0] = 16'hAF6F	;
     642: cos_wave[15:0] = 16'hB010	;
     643: cos_wave[15:0] = 16'hB0B1	;
     644: cos_wave[15:0] = 16'hB153	;
     645: cos_wave[15:0] = 16'hB1F6	;
     646: cos_wave[15:0] = 16'hB29A	;
     647: cos_wave[15:0] = 16'hB33E	;
     648: cos_wave[15:0] = 16'hB3E4	;
     649: cos_wave[15:0] = 16'hB48A	;
     650: cos_wave[15:0] = 16'hB531	;
     651: cos_wave[15:0] = 16'hB5D8	;
     652: cos_wave[15:0] = 16'hB681	;
     653: cos_wave[15:0] = 16'hB72A	;
     654: cos_wave[15:0] = 16'hB7D3	;
     655: cos_wave[15:0] = 16'hB87E	;
     656: cos_wave[15:0] = 16'hB929	;
     657: cos_wave[15:0] = 16'hB9D5	;
     658: cos_wave[15:0] = 16'hBA82	;
     659: cos_wave[15:0] = 16'hBB2F	;
     660: cos_wave[15:0] = 16'hBBDE	;
     661: cos_wave[15:0] = 16'hBC8C	;
     662: cos_wave[15:0] = 16'hBD3C	;
     663: cos_wave[15:0] = 16'hBDEC	;
     664: cos_wave[15:0] = 16'hBE9D	;
     665: cos_wave[15:0] = 16'hBF4E	;
     666: cos_wave[15:0] = 16'hC000	;
     667: cos_wave[15:0] = 16'hC0B3	;
     668: cos_wave[15:0] = 16'hC167	;
     669: cos_wave[15:0] = 16'hC21B	;
     670: cos_wave[15:0] = 16'hC2D0	;
     671: cos_wave[15:0] = 16'hC385	;
     672: cos_wave[15:0] = 16'hC43B	;
     673: cos_wave[15:0] = 16'hC4F1	;
     674: cos_wave[15:0] = 16'hC5A8	;
     675: cos_wave[15:0] = 16'hC660	;
     676: cos_wave[15:0] = 16'hC718	;
     677: cos_wave[15:0] = 16'hC7D1	;
     678: cos_wave[15:0] = 16'hC88B	;
     679: cos_wave[15:0] = 16'hC945	;
     680: cos_wave[15:0] = 16'hC9FF	;
     681: cos_wave[15:0] = 16'hCABB	;
     682: cos_wave[15:0] = 16'hCB76	;
     683: cos_wave[15:0] = 16'hCC32	;
     684: cos_wave[15:0] = 16'hCCEF	;
     685: cos_wave[15:0] = 16'hCDAC	;
     686: cos_wave[15:0] = 16'hCE6A	;
     687: cos_wave[15:0] = 16'hCF28	;
     688: cos_wave[15:0] = 16'hCFE7	;
     689: cos_wave[15:0] = 16'hD0A6	;
     690: cos_wave[15:0] = 16'hD166	;
     691: cos_wave[15:0] = 16'hD226	;
     692: cos_wave[15:0] = 16'hD2E7	;
     693: cos_wave[15:0] = 16'hD3A8	;
     694: cos_wave[15:0] = 16'hD469	;
     695: cos_wave[15:0] = 16'hD52B	;
     696: cos_wave[15:0] = 16'hD5EE	;
     697: cos_wave[15:0] = 16'hD6B1	;
     698: cos_wave[15:0] = 16'hD774	;
     699: cos_wave[15:0] = 16'hD838	;
     700: cos_wave[15:0] = 16'hD8FC	;
     701: cos_wave[15:0] = 16'hD9C0	;
     702: cos_wave[15:0] = 16'hDA85	;
     703: cos_wave[15:0] = 16'hDB4A	;
     704: cos_wave[15:0] = 16'hDC10	;
     705: cos_wave[15:0] = 16'hDCD6	;
     706: cos_wave[15:0] = 16'hDD9C	;
     707: cos_wave[15:0] = 16'hDE63	;
     708: cos_wave[15:0] = 16'hDF2A	;
     709: cos_wave[15:0] = 16'hDFF1	;
     710: cos_wave[15:0] = 16'hE0B9	;
     711: cos_wave[15:0] = 16'hE181	;
     712: cos_wave[15:0] = 16'hE249	;
     713: cos_wave[15:0] = 16'hE312	;
     714: cos_wave[15:0] = 16'hE3DB	;
     715: cos_wave[15:0] = 16'hE4A4	;
     716: cos_wave[15:0] = 16'hE56D	;
     717: cos_wave[15:0] = 16'hE637	;
     718: cos_wave[15:0] = 16'hE701	;
     719: cos_wave[15:0] = 16'hE7CB	;
     720: cos_wave[15:0] = 16'hE896	;
     721: cos_wave[15:0] = 16'hE961	;
     722: cos_wave[15:0] = 16'hEA2C	;
     723: cos_wave[15:0] = 16'hEAF7	;
     724: cos_wave[15:0] = 16'hEBC2	;
     725: cos_wave[15:0] = 16'hEC8E	;
     726: cos_wave[15:0] = 16'hED5A	;
     727: cos_wave[15:0] = 16'hEE26	;
     728: cos_wave[15:0] = 16'hEEF2	;
     729: cos_wave[15:0] = 16'hEFBE	;
     730: cos_wave[15:0] = 16'hF08B	;
     731: cos_wave[15:0] = 16'hF157	;
     732: cos_wave[15:0] = 16'hF224	;
     733: cos_wave[15:0] = 16'hF2F1	;
     734: cos_wave[15:0] = 16'hF3BE	;
     735: cos_wave[15:0] = 16'hF48B	;
     736: cos_wave[15:0] = 16'hF559	;
     737: cos_wave[15:0] = 16'hF626	;
     738: cos_wave[15:0] = 16'hF6F3	;
     739: cos_wave[15:0] = 16'hF7C1	;
     740: cos_wave[15:0] = 16'hF88F	;
     741: cos_wave[15:0] = 16'hF95D	;
     742: cos_wave[15:0] = 16'hFA2A	;
     743: cos_wave[15:0] = 16'hFAF8	;
     744: cos_wave[15:0] = 16'hFBC6	;
     745: cos_wave[15:0] = 16'hFC94	;
     746: cos_wave[15:0] = 16'hFD62	;
     747: cos_wave[15:0] = 16'hFE30	;
     748: cos_wave[15:0] = 16'hFEFE	;
     749: cos_wave[15:0] = 16'hFFCC	;
     750: cos_wave[15:0] = 16'h009B	;
     751: cos_wave[15:0] = 16'h0169	;
     752: cos_wave[15:0] = 16'h0237	;
     753: cos_wave[15:0] = 16'h0305	;
     754: cos_wave[15:0] = 16'h03D3	;
     755: cos_wave[15:0] = 16'h04A1	;
     756: cos_wave[15:0] = 16'h056F	;
     757: cos_wave[15:0] = 16'h063D	;
     758: cos_wave[15:0] = 16'h070A	;
     759: cos_wave[15:0] = 16'h07D8	;
     760: cos_wave[15:0] = 16'h08A6	;
     761: cos_wave[15:0] = 16'h0973	;
     762: cos_wave[15:0] = 16'h0A41	;
     763: cos_wave[15:0] = 16'h0B0E	;
     764: cos_wave[15:0] = 16'h0BDB	;
     765: cos_wave[15:0] = 16'h0CA9	;
     766: cos_wave[15:0] = 16'h0D76	;
     767: cos_wave[15:0] = 16'h0E42	;
     768: cos_wave[15:0] = 16'h0F0F	;
     769: cos_wave[15:0] = 16'h0FDC	;
     770: cos_wave[15:0] = 16'h10A8	;
     771: cos_wave[15:0] = 16'h1174	;
     772: cos_wave[15:0] = 16'h1241	;
     773: cos_wave[15:0] = 16'h130C	;
     774: cos_wave[15:0] = 16'h13D8	;
     775: cos_wave[15:0] = 16'h14A4	;
     776: cos_wave[15:0] = 16'h156F	;
     777: cos_wave[15:0] = 16'h163A	;
     778: cos_wave[15:0] = 16'h1705	;
     779: cos_wave[15:0] = 16'h17CF	;
     780: cos_wave[15:0] = 16'h189A	;
     781: cos_wave[15:0] = 16'h1964	;
     782: cos_wave[15:0] = 16'h1A2E	;
     783: cos_wave[15:0] = 16'h1AF7	;
     784: cos_wave[15:0] = 16'h1BC1	;
     785: cos_wave[15:0] = 16'h1C8A	;
     786: cos_wave[15:0] = 16'h1D52	;
     787: cos_wave[15:0] = 16'h1E1B	;
     788: cos_wave[15:0] = 16'h1EE3	;
     789: cos_wave[15:0] = 16'h1FAB	;
     790: cos_wave[15:0] = 16'h2072	;
     791: cos_wave[15:0] = 16'h213A	;
     792: cos_wave[15:0] = 16'h2200	;
     793: cos_wave[15:0] = 16'h22C7	;
     794: cos_wave[15:0] = 16'h238D	;
     795: cos_wave[15:0] = 16'h2453	;
     796: cos_wave[15:0] = 16'h2518	;
     797: cos_wave[15:0] = 16'h25DD	;
     798: cos_wave[15:0] = 16'h26A2	;
     799: cos_wave[15:0] = 16'h2766	;
     800: cos_wave[15:0] = 16'h282A	;
     801: cos_wave[15:0] = 16'h28EE	;
     802: cos_wave[15:0] = 16'h29B1	;
     803: cos_wave[15:0] = 16'h2A73	;
     804: cos_wave[15:0] = 16'h2B36	;
     805: cos_wave[15:0] = 16'h2BF7	;
     806: cos_wave[15:0] = 16'h2CB9	;
     807: cos_wave[15:0] = 16'h2D7A	;
     808: cos_wave[15:0] = 16'h2E3A	;
     809: cos_wave[15:0] = 16'h2EFA	;
     810: cos_wave[15:0] = 16'h2FB9	;
     811: cos_wave[15:0] = 16'h3078	;
     812: cos_wave[15:0] = 16'h3137	;
     813: cos_wave[15:0] = 16'h31F5	;
     814: cos_wave[15:0] = 16'h32B2	;
     815: cos_wave[15:0] = 16'h336F	;
     816: cos_wave[15:0] = 16'h342C	;
     817: cos_wave[15:0] = 16'h34E8	;
     818: cos_wave[15:0] = 16'h35A3	;
     819: cos_wave[15:0] = 16'h365E	;
     820: cos_wave[15:0] = 16'h3718	;
     821: cos_wave[15:0] = 16'h37D2	;
     822: cos_wave[15:0] = 16'h388B	;
     823: cos_wave[15:0] = 16'h3944	;
     824: cos_wave[15:0] = 16'h39FC	;
     825: cos_wave[15:0] = 16'h3AB3	;
     826: cos_wave[15:0] = 16'h3B6A	;
     827: cos_wave[15:0] = 16'h3C20	;
     828: cos_wave[15:0] = 16'h3CD6	;
     829: cos_wave[15:0] = 16'h3D8B	;
     830: cos_wave[15:0] = 16'h3E3F	;
     831: cos_wave[15:0] = 16'h3EF3	;
     832: cos_wave[15:0] = 16'h3FA6	;
     833: cos_wave[15:0] = 16'h4059	;
     834: cos_wave[15:0] = 16'h410A	;
     835: cos_wave[15:0] = 16'h41BC	;
     836: cos_wave[15:0] = 16'h426C	;
     837: cos_wave[15:0] = 16'h431C	;
     838: cos_wave[15:0] = 16'h43CB	;
     839: cos_wave[15:0] = 16'h447A	;
     840: cos_wave[15:0] = 16'h4527	;
     841: cos_wave[15:0] = 16'h45D4	;
     842: cos_wave[15:0] = 16'h4681	;
     843: cos_wave[15:0] = 16'h472C	;
     844: cos_wave[15:0] = 16'h47D7	;
     845: cos_wave[15:0] = 16'h4882	;
     846: cos_wave[15:0] = 16'h492B	;
     847: cos_wave[15:0] = 16'h49D4	;
     848: cos_wave[15:0] = 16'h4A7C	;
     849: cos_wave[15:0] = 16'h4B23	;
     850: cos_wave[15:0] = 16'h4BC9	;
     851: cos_wave[15:0] = 16'h4C6F	;
     852: cos_wave[15:0] = 16'h4D14	;
     853: cos_wave[15:0] = 16'h4DB8	;
     854: cos_wave[15:0] = 16'h4E5C	;
     855: cos_wave[15:0] = 16'h4EFE	;
     856: cos_wave[15:0] = 16'h4FA0	;
     857: cos_wave[15:0] = 16'h5041	;
     858: cos_wave[15:0] = 16'h50E1	;
     859: cos_wave[15:0] = 16'h5180	;
     860: cos_wave[15:0] = 16'h521F	;
     861: cos_wave[15:0] = 16'h52BC	;
     862: cos_wave[15:0] = 16'h5359	;
     863: cos_wave[15:0] = 16'h53F5	;
     864: cos_wave[15:0] = 16'h5490	;
     865: cos_wave[15:0] = 16'h552B	;
     866: cos_wave[15:0] = 16'h55C4	;
     867: cos_wave[15:0] = 16'h565D	;
     868: cos_wave[15:0] = 16'h56F4	;
     869: cos_wave[15:0] = 16'h578B	;
     870: cos_wave[15:0] = 16'h5821	;
     871: cos_wave[15:0] = 16'h58B6	;
     872: cos_wave[15:0] = 16'h594A	;
     873: cos_wave[15:0] = 16'h59DD	;
     874: cos_wave[15:0] = 16'h5A70	;
     875: cos_wave[15:0] = 16'h5B01	;
     876: cos_wave[15:0] = 16'h5B91	;
     877: cos_wave[15:0] = 16'h5C21	;
     878: cos_wave[15:0] = 16'h5CB0	;
     879: cos_wave[15:0] = 16'h5D3D	;
     880: cos_wave[15:0] = 16'h5DCA	;
     881: cos_wave[15:0] = 16'h5E56	;
     882: cos_wave[15:0] = 16'h5EE0	;
     883: cos_wave[15:0] = 16'h5F6A	;
     884: cos_wave[15:0] = 16'h5FF3	;
     885: cos_wave[15:0] = 16'h607B	;
     886: cos_wave[15:0] = 16'h6102	;
     887: cos_wave[15:0] = 16'h6188	;
     888: cos_wave[15:0] = 16'h620D	;
     889: cos_wave[15:0] = 16'h6291	;
     890: cos_wave[15:0] = 16'h6314	;
     891: cos_wave[15:0] = 16'h6396	;
     892: cos_wave[15:0] = 16'h6417	;
     893: cos_wave[15:0] = 16'h6497	;
     894: cos_wave[15:0] = 16'h6516	;
     895: cos_wave[15:0] = 16'h6594	;
     896: cos_wave[15:0] = 16'h6611	;
     897: cos_wave[15:0] = 16'h668C	;
     898: cos_wave[15:0] = 16'h6707	;
     899: cos_wave[15:0] = 16'h6781	;
     900: cos_wave[15:0] = 16'h67FA	;
     901: cos_wave[15:0] = 16'h6871	;
     902: cos_wave[15:0] = 16'h68E8	;
     903: cos_wave[15:0] = 16'h695D	;
     904: cos_wave[15:0] = 16'h69D2	;
     905: cos_wave[15:0] = 16'h6A45	;
     906: cos_wave[15:0] = 16'h6AB8	;
     907: cos_wave[15:0] = 16'h6B29	;
     908: cos_wave[15:0] = 16'h6B99	;
     909: cos_wave[15:0] = 16'h6C08	;
     910: cos_wave[15:0] = 16'h6C76	;
     911: cos_wave[15:0] = 16'h6CE3	;
     912: cos_wave[15:0] = 16'h6D4F	;
     913: cos_wave[15:0] = 16'h6DB9	;
     914: cos_wave[15:0] = 16'h6E23	;
     915: cos_wave[15:0] = 16'h6E8B	;
     916: cos_wave[15:0] = 16'h6EF3	;
     917: cos_wave[15:0] = 16'h6F59	;
     918: cos_wave[15:0] = 16'h6FBE	;
     919: cos_wave[15:0] = 16'h7022	;
     920: cos_wave[15:0] = 16'h7085	;
     921: cos_wave[15:0] = 16'h70E6	;
     922: cos_wave[15:0] = 16'h7147	;
     923: cos_wave[15:0] = 16'h71A6	;
     924: cos_wave[15:0] = 16'h7205	;
     925: cos_wave[15:0] = 16'h7262	;
     926: cos_wave[15:0] = 16'h72BE	;
     927: cos_wave[15:0] = 16'h7318	;
     928: cos_wave[15:0] = 16'h7372	;
     929: cos_wave[15:0] = 16'h73CA	;
     930: cos_wave[15:0] = 16'h7422	;
     931: cos_wave[15:0] = 16'h7478	;
     932: cos_wave[15:0] = 16'h74CD	;
     933: cos_wave[15:0] = 16'h7520	;
     934: cos_wave[15:0] = 16'h7573	;
     935: cos_wave[15:0] = 16'h75C4	;
     936: cos_wave[15:0] = 16'h7614	;
     937: cos_wave[15:0] = 16'h7663	;
     938: cos_wave[15:0] = 16'h76B1	;
     939: cos_wave[15:0] = 16'h76FD	;
     940: cos_wave[15:0] = 16'h7749	;
     941: cos_wave[15:0] = 16'h7793	;
     942: cos_wave[15:0] = 16'h77DC	;
     943: cos_wave[15:0] = 16'h7824	;
     944: cos_wave[15:0] = 16'h786A	;
     945: cos_wave[15:0] = 16'h78AF	;
     946: cos_wave[15:0] = 16'h78F3	;
     947: cos_wave[15:0] = 16'h7936	;
     948: cos_wave[15:0] = 16'h7978	;
     949: cos_wave[15:0] = 16'h79B8	;
     950: cos_wave[15:0] = 16'h79F7	;
     951: cos_wave[15:0] = 16'h7A35	;
     952: cos_wave[15:0] = 16'h7A72	;
     953: cos_wave[15:0] = 16'h7AAD	;
     954: cos_wave[15:0] = 16'h7AE7	;
     955: cos_wave[15:0] = 16'h7B20	;
     956: cos_wave[15:0] = 16'h7B58	;
     957: cos_wave[15:0] = 16'h7B8E	;
     958: cos_wave[15:0] = 16'h7BC4	;
     959: cos_wave[15:0] = 16'h7BF8	;
     960: cos_wave[15:0] = 16'h7C2A	;
     961: cos_wave[15:0] = 16'h7C5C	;
     962: cos_wave[15:0] = 16'h7C8C	;
     963: cos_wave[15:0] = 16'h7CBB	;
     964: cos_wave[15:0] = 16'h7CE8	;
     965: cos_wave[15:0] = 16'h7D15	;
     966: cos_wave[15:0] = 16'h7D40	;
     967: cos_wave[15:0] = 16'h7D6A	;
     968: cos_wave[15:0] = 16'h7D92	;
     969: cos_wave[15:0] = 16'h7DB9	;
     970: cos_wave[15:0] = 16'h7DDF	;
     971: cos_wave[15:0] = 16'h7E04	;
     972: cos_wave[15:0] = 16'h7E28	;
     973: cos_wave[15:0] = 16'h7E4A	;
     974: cos_wave[15:0] = 16'h7E6B	;
     975: cos_wave[15:0] = 16'h7E8A	;
     976: cos_wave[15:0] = 16'h7EA9	;
     977: cos_wave[15:0] = 16'h7EC6	;
     978: cos_wave[15:0] = 16'h7EE2	;
     979: cos_wave[15:0] = 16'h7EFC	;
     980: cos_wave[15:0] = 16'h7F15	;
     981: cos_wave[15:0] = 16'h7F2D	;
     982: cos_wave[15:0] = 16'h7F44	;
     983: cos_wave[15:0] = 16'h7F59	;
     984: cos_wave[15:0] = 16'h7F6D	;
     985: cos_wave[15:0] = 16'h7F80	;
     986: cos_wave[15:0] = 16'h7F92	;
     987: cos_wave[15:0] = 16'h7FA2	;
     988: cos_wave[15:0] = 16'h7FB1	;
     989: cos_wave[15:0] = 16'h7FBE	;
     990: cos_wave[15:0] = 16'h7FCB	;
     991: cos_wave[15:0] = 16'h7FD6	;
     992: cos_wave[15:0] = 16'h7FDF	;
     993: cos_wave[15:0] = 16'h7FE8	;
     994: cos_wave[15:0] = 16'h7FEF	;
     995: cos_wave[15:0] = 16'h7FF5	;
     996: cos_wave[15:0] = 16'h7FF9	;
     997: cos_wave[15:0] = 16'h7FFC	;
     998: cos_wave[15:0] = 16'h7FFE	;
     999: cos_wave[15:0] = 16'h7FFF	;
     endcase
end
//    
endmodule
