module pure_sin_table(
     input              sclk,
     input              rst_n,
     output wire [15:0] pure_sin
    );
//
assign pure_sin[15:0] = sin_wave[15:0];
//
parameter lim = 999;
//
reg  [9:0] cnt;
reg [15:0] sin_wave;
//
always @(posedge sclk or negedge rst_n)
begin
     if (!rst_n)        cnt <= 0 ;
     else if (lim==cnt) cnt <= 0 ;
     else               cnt <= cnt+1 ; 
end
//
always @(posedge sclk or negedge rst_n)
begin
     if (!rst_n) sin_wave[15:0] = 16'h0000 ;
     else
     case(cnt)
     0	: sin_wave[15:0] = 16'h0000	;
     1	: sin_wave[15:0] = 16'h00CE	;
     2	: sin_wave[15:0] = 16'h019C	;
     3	: sin_wave[15:0] = 16'h026A	;
     4	: sin_wave[15:0] = 16'h0338	;
     5	: sin_wave[15:0] = 16'h0406	;
     6	: sin_wave[15:0] = 16'h04D4	;
     7	: sin_wave[15:0] = 16'h05A2	;
     8	: sin_wave[15:0] = 16'h0670	;
     9	: sin_wave[15:0] = 16'h073E	;
     10	: sin_wave[15:0] = 16'h080C	;
     11	: sin_wave[15:0] = 16'h08D9	;
     12	: sin_wave[15:0] = 16'h09A7	;
     13	: sin_wave[15:0] = 16'h0A74	;
     14	: sin_wave[15:0] = 16'h0B41	;
     15	: sin_wave[15:0] = 16'h0C0F	;
     16	: sin_wave[15:0] = 16'h0CDC	;
     17	: sin_wave[15:0] = 16'h0DA9	;
     18	: sin_wave[15:0] = 16'h0E76	;
     19	: sin_wave[15:0] = 16'h0F42	;
     20	: sin_wave[15:0] = 16'h100F	;
     21	: sin_wave[15:0] = 16'h10DB	;
     22	: sin_wave[15:0] = 16'h11A7	;
     23	: sin_wave[15:0] = 16'h1273	;
     24	: sin_wave[15:0] = 16'h133F	;
     25	: sin_wave[15:0] = 16'h140B	;
     26	: sin_wave[15:0] = 16'h14D6	;
     27	: sin_wave[15:0] = 16'h15A2	;
     28	: sin_wave[15:0] = 16'h166D	;
     29	: sin_wave[15:0] = 16'h1737	;
     30	: sin_wave[15:0] = 16'h1802	;
     31	: sin_wave[15:0] = 16'h18CC	;
     32	: sin_wave[15:0] = 16'h1996	;
     33	: sin_wave[15:0] = 16'h1A60	;
     34	: sin_wave[15:0] = 16'h1B2A	;
     35	: sin_wave[15:0] = 16'h1BF3	;
     36	: sin_wave[15:0] = 16'h1CBC	;
     37	: sin_wave[15:0] = 16'h1D85	;
     38	: sin_wave[15:0] = 16'h1E4D	;
     39	: sin_wave[15:0] = 16'h1F15	;
     40	: sin_wave[15:0] = 16'h1FDD	;
     41	: sin_wave[15:0] = 16'h20A4	;
     42	: sin_wave[15:0] = 16'h216B	;
     43	: sin_wave[15:0] = 16'h2232	;
     44	: sin_wave[15:0] = 16'h22F9	;
     45	: sin_wave[15:0] = 16'h23BF	;
     46	: sin_wave[15:0] = 16'h2484	;
     47	: sin_wave[15:0] = 16'h254A	;
     48	: sin_wave[15:0] = 16'h260F	;
     49	: sin_wave[15:0] = 16'h26D3	;
     50	: sin_wave[15:0] = 16'h2797	;
     51	: sin_wave[15:0] = 16'h285B	;
     52	: sin_wave[15:0] = 16'h291F	;
     53	: sin_wave[15:0] = 16'h29E1	;
     54	: sin_wave[15:0] = 16'h2AA4	;
     55	: sin_wave[15:0] = 16'h2B66	;
     56	: sin_wave[15:0] = 16'h2C28	;
     57	: sin_wave[15:0] = 16'h2CE9	;
     58	: sin_wave[15:0] = 16'h2DAA	;
     59	: sin_wave[15:0] = 16'h2E6A	;
     60	: sin_wave[15:0] = 16'h2F2A	;
     61	: sin_wave[15:0] = 16'h2FE9	;
     62	: sin_wave[15:0] = 16'h30A8	;
     63	: sin_wave[15:0] = 16'h3166	;
     64	: sin_wave[15:0] = 16'h3224	;
     65	: sin_wave[15:0] = 16'h32E2	;
     66	: sin_wave[15:0] = 16'h339E	;
     67	: sin_wave[15:0] = 16'h345B	;
     68	: sin_wave[15:0] = 16'h3517	;
     69	: sin_wave[15:0] = 16'h35D2	;
     70	: sin_wave[15:0] = 16'h368D	;
     71	: sin_wave[15:0] = 16'h3747	;
     72	: sin_wave[15:0] = 16'h3800	;
     73	: sin_wave[15:0] = 16'h38B9	;
     74	: sin_wave[15:0] = 16'h3972	;
     75	: sin_wave[15:0] = 16'h3A2A	;
     76	: sin_wave[15:0] = 16'h3AE1	;
     77	: sin_wave[15:0] = 16'h3B98	;
     78	: sin_wave[15:0] = 16'h3C4E	;
     79	: sin_wave[15:0] = 16'h3D03	;
     80	: sin_wave[15:0] = 16'h3DB8	;
     81	: sin_wave[15:0] = 16'h3E6C	;
     82	: sin_wave[15:0] = 16'h3F20	;
     83	: sin_wave[15:0] = 16'h3FD3	;
     84	: sin_wave[15:0] = 16'h4085	;
     85	: sin_wave[15:0] = 16'h4137	;
     86	: sin_wave[15:0] = 16'h41E8	;
     87	: sin_wave[15:0] = 16'h4298	;
     88	: sin_wave[15:0] = 16'h4348	;
     89	: sin_wave[15:0] = 16'h43F7	;
     90	: sin_wave[15:0] = 16'h44A5	;
     91	: sin_wave[15:0] = 16'h4553	;
     92	: sin_wave[15:0] = 16'h4600	;
     93	: sin_wave[15:0] = 16'h46AC	;
     94	: sin_wave[15:0] = 16'h4757	;
     95	: sin_wave[15:0] = 16'h4802	;
     96	: sin_wave[15:0] = 16'h48AC	;
     97	: sin_wave[15:0] = 16'h4955	;
     98	: sin_wave[15:0] = 16'h49FE	;
     99	: sin_wave[15:0] = 16'h4AA6	;
     100: sin_wave[15:0] = 16'h4B4D	;
     101: sin_wave[15:0] = 16'h4BF3	;
     102: sin_wave[15:0] = 16'h4C98	;
     103: sin_wave[15:0] = 16'h4D3D	;
     104: sin_wave[15:0] = 16'h4DE1	;
     105: sin_wave[15:0] = 16'h4E84	;
     106: sin_wave[15:0] = 16'h4F27	;
     107: sin_wave[15:0] = 16'h4FC8	;
     108: sin_wave[15:0] = 16'h5069	;
     109: sin_wave[15:0] = 16'h5109	;
     110: sin_wave[15:0] = 16'h51A8	;
     111: sin_wave[15:0] = 16'h5246	;
     112: sin_wave[15:0] = 16'h52E4	;
     113: sin_wave[15:0] = 16'h5380	;
     114: sin_wave[15:0] = 16'h541C	;
     115: sin_wave[15:0] = 16'h54B7	;
     116: sin_wave[15:0] = 16'h5551	;
     117: sin_wave[15:0] = 16'h55EA	;
     118: sin_wave[15:0] = 16'h5683	;
     119: sin_wave[15:0] = 16'h571A	;
     120: sin_wave[15:0] = 16'h57B1	;
     121: sin_wave[15:0] = 16'h5846	;
     122: sin_wave[15:0] = 16'h58DB	;
     123: sin_wave[15:0] = 16'h596F	;
     124: sin_wave[15:0] = 16'h5A02	;
     125: sin_wave[15:0] = 16'h5A94	;
     126: sin_wave[15:0] = 16'h5B25	;
     127: sin_wave[15:0] = 16'h5BB5	;
     128: sin_wave[15:0] = 16'h5C45	;
     129: sin_wave[15:0] = 16'h5CD3	;
     130: sin_wave[15:0] = 16'h5D60	;
     131: sin_wave[15:0] = 16'h5DED	;
     132: sin_wave[15:0] = 16'h5E78	;
     133: sin_wave[15:0] = 16'h5F03	;
     134: sin_wave[15:0] = 16'h5F8D	;
     135: sin_wave[15:0] = 16'h6015	;
     136: sin_wave[15:0] = 16'h609D	;
     137: sin_wave[15:0] = 16'h6124	;
     138: sin_wave[15:0] = 16'h61A9	;
     139: sin_wave[15:0] = 16'h622E	;
     140: sin_wave[15:0] = 16'h62B2	;
     141: sin_wave[15:0] = 16'h6335	;
     142: sin_wave[15:0] = 16'h63B6	;
     143: sin_wave[15:0] = 16'h6437	;
     144: sin_wave[15:0] = 16'h64B7	;
     145: sin_wave[15:0] = 16'h6535	;
     146: sin_wave[15:0] = 16'h65B3	;
     147: sin_wave[15:0] = 16'h6630	;
     148: sin_wave[15:0] = 16'h66AB	;
     149: sin_wave[15:0] = 16'h6726	;
     150: sin_wave[15:0] = 16'h679F	;
     151: sin_wave[15:0] = 16'h6818	;
     152: sin_wave[15:0] = 16'h688F	;
     153: sin_wave[15:0] = 16'h6905	;
     154: sin_wave[15:0] = 16'h697B	;
     155: sin_wave[15:0] = 16'h69EF	;
     156: sin_wave[15:0] = 16'h6A62	;
     157: sin_wave[15:0] = 16'h6AD4	;
     158: sin_wave[15:0] = 16'h6B45	;
     159: sin_wave[15:0] = 16'h6BB5	;
     160: sin_wave[15:0] = 16'h6C24	;
     161: sin_wave[15:0] = 16'h6C91	;
     162: sin_wave[15:0] = 16'h6CFE	;
     163: sin_wave[15:0] = 16'h6D6A	;
     164: sin_wave[15:0] = 16'h6DD4	;
     165: sin_wave[15:0] = 16'h6E3D	;
     166: sin_wave[15:0] = 16'h6EA5	;
     167: sin_wave[15:0] = 16'h6F0C	;
     168: sin_wave[15:0] = 16'h6F72	;
     169: sin_wave[15:0] = 16'h6FD7	;
     170: sin_wave[15:0] = 16'h703B	;
     171: sin_wave[15:0] = 16'h709D	;
     172: sin_wave[15:0] = 16'h70FF	;
     173: sin_wave[15:0] = 16'h715F	;
     174: sin_wave[15:0] = 16'h71BE	;
     175: sin_wave[15:0] = 16'h721C	;
     176: sin_wave[15:0] = 16'h7279	;
     177: sin_wave[15:0] = 16'h72D4	;
     178: sin_wave[15:0] = 16'h732F	;
     179: sin_wave[15:0] = 16'h7388	;
     180: sin_wave[15:0] = 16'h73E0	;
     181: sin_wave[15:0] = 16'h7437	;
     182: sin_wave[15:0] = 16'h748D	;
     183: sin_wave[15:0] = 16'h74E2	;
     184: sin_wave[15:0] = 16'h7535	;
     185: sin_wave[15:0] = 16'h7587	;
     186: sin_wave[15:0] = 16'h75D8	;
     187: sin_wave[15:0] = 16'h7628	;
     188: sin_wave[15:0] = 16'h7677	;
     189: sin_wave[15:0] = 16'h76C4	;
     190: sin_wave[15:0] = 16'h7710	;
     191: sin_wave[15:0] = 16'h775B	;
     192: sin_wave[15:0] = 16'h77A5	;
     193: sin_wave[15:0] = 16'h77EE	;
     194: sin_wave[15:0] = 16'h7835	;
     195: sin_wave[15:0] = 16'h787B	;
     196: sin_wave[15:0] = 16'h78C0	;
     197: sin_wave[15:0] = 16'h7904	;
     198: sin_wave[15:0] = 16'h7947	;
     199: sin_wave[15:0] = 16'h7988	;
     200: sin_wave[15:0] = 16'h79C8	;
     201: sin_wave[15:0] = 16'h7A07	;
     202: sin_wave[15:0] = 16'h7A44	;
     203: sin_wave[15:0] = 16'h7A81	;
     204: sin_wave[15:0] = 16'h7ABC	;
     205: sin_wave[15:0] = 16'h7AF6	;
     206: sin_wave[15:0] = 16'h7B2E	;
     207: sin_wave[15:0] = 16'h7B66	;
     208: sin_wave[15:0] = 16'h7B9C	;
     209: sin_wave[15:0] = 16'h7BD1	;
     210: sin_wave[15:0] = 16'h7C04	;
     211: sin_wave[15:0] = 16'h7C37	;
     212: sin_wave[15:0] = 16'h7C68	;
     213: sin_wave[15:0] = 16'h7C98	;
     214: sin_wave[15:0] = 16'h7CC6	;
     215: sin_wave[15:0] = 16'h7CF4	;
     216: sin_wave[15:0] = 16'h7D20	;
     217: sin_wave[15:0] = 16'h7D4A	;
     218: sin_wave[15:0] = 16'h7D74	;
     219: sin_wave[15:0] = 16'h7D9C	;
     220: sin_wave[15:0] = 16'h7DC3	;
     221: sin_wave[15:0] = 16'h7DE9	;
     222: sin_wave[15:0] = 16'h7E0D	;
     223: sin_wave[15:0] = 16'h7E30	;
     224: sin_wave[15:0] = 16'h7E52	;
     225: sin_wave[15:0] = 16'h7E73	;
     226: sin_wave[15:0] = 16'h7E92	;
     227: sin_wave[15:0] = 16'h7EB0	;
     228: sin_wave[15:0] = 16'h7ECD	;
     229: sin_wave[15:0] = 16'h7EE8	;
     230: sin_wave[15:0] = 16'h7F03	;
     231: sin_wave[15:0] = 16'h7F1B	;
     232: sin_wave[15:0] = 16'h7F33	;
     233: sin_wave[15:0] = 16'h7F49	;
     234: sin_wave[15:0] = 16'h7F5E	;
     235: sin_wave[15:0] = 16'h7F72	;
     236: sin_wave[15:0] = 16'h7F85	;
     237: sin_wave[15:0] = 16'h7F96	;
     238: sin_wave[15:0] = 16'h7FA6	;
     239: sin_wave[15:0] = 16'h7FB4	;
     240: sin_wave[15:0] = 16'h7FC1	;
     241: sin_wave[15:0] = 16'h7FCD	;
     242: sin_wave[15:0] = 16'h7FD8	;
     243: sin_wave[15:0] = 16'h7FE1	;
     244: sin_wave[15:0] = 16'h7FEA	;
     245: sin_wave[15:0] = 16'h7FF0	;
     246: sin_wave[15:0] = 16'h7FF6	;
     247: sin_wave[15:0] = 16'h7FFA	;
     248: sin_wave[15:0] = 16'h7FFD	;
     249: sin_wave[15:0] = 16'h7FFF	;
     250: sin_wave[15:0] = 16'h7FFF	;
     251: sin_wave[15:0] = 16'h7FFE	;
     252: sin_wave[15:0] = 16'h7FFC	;
     253: sin_wave[15:0] = 16'h7FF8	;
     254: sin_wave[15:0] = 16'h7FF3	;
     255: sin_wave[15:0] = 16'h7FED	;
     256: sin_wave[15:0] = 16'h7FE6	;
     257: sin_wave[15:0] = 16'h7FDD	;
     258: sin_wave[15:0] = 16'h7FD3	;
     259: sin_wave[15:0] = 16'h7FC8	;
     260: sin_wave[15:0] = 16'h7FBB	;
     261: sin_wave[15:0] = 16'h7FAD	;
     262: sin_wave[15:0] = 16'h7F9E	;
     263: sin_wave[15:0] = 16'h7F8D	;
     264: sin_wave[15:0] = 16'h7F7B	;
     265: sin_wave[15:0] = 16'h7F68	;
     266: sin_wave[15:0] = 16'h7F54	;
     267: sin_wave[15:0] = 16'h7F3E	;
     268: sin_wave[15:0] = 16'h7F27	;
     269: sin_wave[15:0] = 16'h7F0F	;
     270: sin_wave[15:0] = 16'h7EF6	;
     271: sin_wave[15:0] = 16'h7EDB	;
     272: sin_wave[15:0] = 16'h7EBF	;
     273: sin_wave[15:0] = 16'h7EA1	;
     274: sin_wave[15:0] = 16'h7E83	;
     275: sin_wave[15:0] = 16'h7E63	;
     276: sin_wave[15:0] = 16'h7E41	;
     277: sin_wave[15:0] = 16'h7E1F	;
     278: sin_wave[15:0] = 16'h7DFB	;
     279: sin_wave[15:0] = 16'h7DD6	;
     280: sin_wave[15:0] = 16'h7DB0	;
     281: sin_wave[15:0] = 16'h7D88	;
     282: sin_wave[15:0] = 16'h7D5F	;
     283: sin_wave[15:0] = 16'h7D35	;
     284: sin_wave[15:0] = 16'h7D0A	;
     285: sin_wave[15:0] = 16'h7CDD	;
     286: sin_wave[15:0] = 16'h7CAF	;
     287: sin_wave[15:0] = 16'h7C80	;
     288: sin_wave[15:0] = 16'h7C4F	;
     289: sin_wave[15:0] = 16'h7C1E	;
     290: sin_wave[15:0] = 16'h7BEB	;
     291: sin_wave[15:0] = 16'h7BB6	;
     292: sin_wave[15:0] = 16'h7B81	;
     293: sin_wave[15:0] = 16'h7B4A	;
     294: sin_wave[15:0] = 16'h7B12	;
     295: sin_wave[15:0] = 16'h7AD9	;
     296: sin_wave[15:0] = 16'h7A9E	;
     297: sin_wave[15:0] = 16'h7A63	;
     298: sin_wave[15:0] = 16'h7A26	;
     299: sin_wave[15:0] = 16'h79E8	;
     300: sin_wave[15:0] = 16'h79A8	;
     301: sin_wave[15:0] = 16'h7967	;
     302: sin_wave[15:0] = 16'h7926	;
     303: sin_wave[15:0] = 16'h78E2	;
     304: sin_wave[15:0] = 16'h789E	;
     305: sin_wave[15:0] = 16'h7858	;
     306: sin_wave[15:0] = 16'h7812	;
     307: sin_wave[15:0] = 16'h77CA	;
     308: sin_wave[15:0] = 16'h7780	;
     309: sin_wave[15:0] = 16'h7736	;
     310: sin_wave[15:0] = 16'h76EA	;
     311: sin_wave[15:0] = 16'h769E	;
     312: sin_wave[15:0] = 16'h7650	;
     313: sin_wave[15:0] = 16'h7600	;
     314: sin_wave[15:0] = 16'h75B0	;
     315: sin_wave[15:0] = 16'h755E	;
     316: sin_wave[15:0] = 16'h750B	;
     317: sin_wave[15:0] = 16'h74B7	;
     318: sin_wave[15:0] = 16'h7462	;
     319: sin_wave[15:0] = 16'h740C	;
     320: sin_wave[15:0] = 16'h73B4	;
     321: sin_wave[15:0] = 16'h735C	;
     322: sin_wave[15:0] = 16'h7302	;
     323: sin_wave[15:0] = 16'h72A7	;
     324: sin_wave[15:0] = 16'h724B	;
     325: sin_wave[15:0] = 16'h71ED	;
     326: sin_wave[15:0] = 16'h718F	;
     327: sin_wave[15:0] = 16'h712F	;
     328: sin_wave[15:0] = 16'h70CE	;
     329: sin_wave[15:0] = 16'h706C	;
     330: sin_wave[15:0] = 16'h7009	;
     331: sin_wave[15:0] = 16'h6FA5	;
     332: sin_wave[15:0] = 16'h6F40	;
     333: sin_wave[15:0] = 16'h6ED9	;
     334: sin_wave[15:0] = 16'h6E71	;
     335: sin_wave[15:0] = 16'h6E09	;
     336: sin_wave[15:0] = 16'h6D9F	;
     337: sin_wave[15:0] = 16'h6D34	;
     338: sin_wave[15:0] = 16'h6CC8	;
     339: sin_wave[15:0] = 16'h6C5B	;
     340: sin_wave[15:0] = 16'h6BEC	;
     341: sin_wave[15:0] = 16'h6B7D	;
     342: sin_wave[15:0] = 16'h6B0D	;
     343: sin_wave[15:0] = 16'h6A9B	;
     344: sin_wave[15:0] = 16'h6A29	;
     345: sin_wave[15:0] = 16'h69B5	;
     346: sin_wave[15:0] = 16'h6940	;
     347: sin_wave[15:0] = 16'h68CA	;
     348: sin_wave[15:0] = 16'h6854	;
     349: sin_wave[15:0] = 16'h67DC	;
     350: sin_wave[15:0] = 16'h6763	;
     351: sin_wave[15:0] = 16'h66E9	;
     352: sin_wave[15:0] = 16'h666E	;
     353: sin_wave[15:0] = 16'h65F1	;
     354: sin_wave[15:0] = 16'h6574	;
     355: sin_wave[15:0] = 16'h64F6	;
     356: sin_wave[15:0] = 16'h6477	;
     357: sin_wave[15:0] = 16'h63F7	;
     358: sin_wave[15:0] = 16'h6375	;
     359: sin_wave[15:0] = 16'h62F3	;
     360: sin_wave[15:0] = 16'h6270	;
     361: sin_wave[15:0] = 16'h61EC	;
     362: sin_wave[15:0] = 16'h6167	;
     363: sin_wave[15:0] = 16'h60E0	;
     364: sin_wave[15:0] = 16'h6059	;
     365: sin_wave[15:0] = 16'h5FD1	;
     366: sin_wave[15:0] = 16'h5F48	;
     367: sin_wave[15:0] = 16'h5EBE	;
     368: sin_wave[15:0] = 16'h5E33	;
     369: sin_wave[15:0] = 16'h5DA7	;
     370: sin_wave[15:0] = 16'h5D1A	;
     371: sin_wave[15:0] = 16'h5C8C	;
     372: sin_wave[15:0] = 16'h5BFD	;
     373: sin_wave[15:0] = 16'h5B6D	;
     374: sin_wave[15:0] = 16'h5ADD	;
     375: sin_wave[15:0] = 16'h5A4B	;
     376: sin_wave[15:0] = 16'h59B9	;
     377: sin_wave[15:0] = 16'h5925	;
     378: sin_wave[15:0] = 16'h5891	;
     379: sin_wave[15:0] = 16'h57FC	;
     380: sin_wave[15:0] = 16'h5765	;
     381: sin_wave[15:0] = 16'h56CE	;
     382: sin_wave[15:0] = 16'h5637	;
     383: sin_wave[15:0] = 16'h559E	;
     384: sin_wave[15:0] = 16'h5504	;
     385: sin_wave[15:0] = 16'h546A	;
     386: sin_wave[15:0] = 16'h53CE	;
     387: sin_wave[15:0] = 16'h5332	;
     388: sin_wave[15:0] = 16'h5295	;
     389: sin_wave[15:0] = 16'h51F7	;
     390: sin_wave[15:0] = 16'h5158	;
     391: sin_wave[15:0] = 16'h50B9	;
     392: sin_wave[15:0] = 16'h5019	;
     393: sin_wave[15:0] = 16'h4F77	;
     394: sin_wave[15:0] = 16'h4ED5	;
     395: sin_wave[15:0] = 16'h4E33	;
     396: sin_wave[15:0] = 16'h4D8F	;
     397: sin_wave[15:0] = 16'h4CEB	;
     398: sin_wave[15:0] = 16'h4C46	;
     399: sin_wave[15:0] = 16'h4BA0	;
     400: sin_wave[15:0] = 16'h4AF9	;
     401: sin_wave[15:0] = 16'h4A52	;
     402: sin_wave[15:0] = 16'h49AA	;
     403: sin_wave[15:0] = 16'h4901	;
     404: sin_wave[15:0] = 16'h4857	;
     405: sin_wave[15:0] = 16'h47AD	;
     406: sin_wave[15:0] = 16'h4702	;
     407: sin_wave[15:0] = 16'h4656	;
     408: sin_wave[15:0] = 16'h45A9	;
     409: sin_wave[15:0] = 16'h44FC	;
     410: sin_wave[15:0] = 16'h444E	;
     411: sin_wave[15:0] = 16'h439F	;
     412: sin_wave[15:0] = 16'h42F0	;
     413: sin_wave[15:0] = 16'h4240	;
     414: sin_wave[15:0] = 16'h418F	;
     415: sin_wave[15:0] = 16'h40DE	;
     416: sin_wave[15:0] = 16'h402C	;
     417: sin_wave[15:0] = 16'h3F79	;
     418: sin_wave[15:0] = 16'h3EC6	;
     419: sin_wave[15:0] = 16'h3E12	;
     420: sin_wave[15:0] = 16'h3D5E	;
     421: sin_wave[15:0] = 16'h3CA9	;
     422: sin_wave[15:0] = 16'h3BF3	;
     423: sin_wave[15:0] = 16'h3B3C	;
     424: sin_wave[15:0] = 16'h3A85	;
     425: sin_wave[15:0] = 16'h39CE	;
     426: sin_wave[15:0] = 16'h3916	;
     427: sin_wave[15:0] = 16'h385D	;
     428: sin_wave[15:0] = 16'h37A4	;
     429: sin_wave[15:0] = 16'h36EA	;
     430: sin_wave[15:0] = 16'h362F	;
     431: sin_wave[15:0] = 16'h3574	;
     432: sin_wave[15:0] = 16'h34B9	;
     433: sin_wave[15:0] = 16'h33FD	;
     434: sin_wave[15:0] = 16'h3340	;
     435: sin_wave[15:0] = 16'h3283	;
     436: sin_wave[15:0] = 16'h31C5	;
     437: sin_wave[15:0] = 16'h3107	;
     438: sin_wave[15:0] = 16'h3049	;
     439: sin_wave[15:0] = 16'h2F8A	;
     440: sin_wave[15:0] = 16'h2ECA	;
     441: sin_wave[15:0] = 16'h2E0A	;
     442: sin_wave[15:0] = 16'h2D49	;
     443: sin_wave[15:0] = 16'h2C88	;
     444: sin_wave[15:0] = 16'h2BC7	;
     445: sin_wave[15:0] = 16'h2B05	;
     446: sin_wave[15:0] = 16'h2A43	;
     447: sin_wave[15:0] = 16'h2980	;
     448: sin_wave[15:0] = 16'h28BD	;
     449: sin_wave[15:0] = 16'h27F9	;
     450: sin_wave[15:0] = 16'h2735	;
     451: sin_wave[15:0] = 16'h2671	;
     452: sin_wave[15:0] = 16'h25AC	;
     453: sin_wave[15:0] = 16'h24E7	;
     454: sin_wave[15:0] = 16'h2422	;
     455: sin_wave[15:0] = 16'h235C	;
     456: sin_wave[15:0] = 16'h2295	;
     457: sin_wave[15:0] = 16'h21CF	;
     458: sin_wave[15:0] = 16'h2108	;
     459: sin_wave[15:0] = 16'h2041	;
     460: sin_wave[15:0] = 16'h1F79	;
     461: sin_wave[15:0] = 16'h1EB1	;
     462: sin_wave[15:0] = 16'h1DE9	;
     463: sin_wave[15:0] = 16'h1D20	;
     464: sin_wave[15:0] = 16'h1C57	;
     465: sin_wave[15:0] = 16'h1B8E	;
     466: sin_wave[15:0] = 16'h1AC5	;
     467: sin_wave[15:0] = 16'h19FB	;
     468: sin_wave[15:0] = 16'h1931	;
     469: sin_wave[15:0] = 16'h1867	;
     470: sin_wave[15:0] = 16'h179D	;
     471: sin_wave[15:0] = 16'h16D2	;
     472: sin_wave[15:0] = 16'h1607	;
     473: sin_wave[15:0] = 16'h153C	;
     474: sin_wave[15:0] = 16'h1471	;
     475: sin_wave[15:0] = 16'h13A5	;
     476: sin_wave[15:0] = 16'h12D9	;
     477: sin_wave[15:0] = 16'h120E	;
     478: sin_wave[15:0] = 16'h1141	;
     479: sin_wave[15:0] = 16'h1075	;
     480: sin_wave[15:0] = 16'h0FA9	;
     481: sin_wave[15:0] = 16'h0EDC	;
     482: sin_wave[15:0] = 16'h0E0F	;
     483: sin_wave[15:0] = 16'h0D42	;
     484: sin_wave[15:0] = 16'h0C75	;
     485: sin_wave[15:0] = 16'h0BA8	;
     486: sin_wave[15:0] = 16'h0ADB	;
     487: sin_wave[15:0] = 16'h0A0D	;
     488: sin_wave[15:0] = 16'h0940	;
     489: sin_wave[15:0] = 16'h0872	;
     490: sin_wave[15:0] = 16'h07A5	;
     491: sin_wave[15:0] = 16'h06D7	;
     492: sin_wave[15:0] = 16'h0609	;
     493: sin_wave[15:0] = 16'h053B	;
     494: sin_wave[15:0] = 16'h046D	;
     495: sin_wave[15:0] = 16'h039F	;
     496: sin_wave[15:0] = 16'h02D1	;
     497: sin_wave[15:0] = 16'h0203	;
     498: sin_wave[15:0] = 16'h0135	;
     499: sin_wave[15:0] = 16'h0067	;
     500: sin_wave[15:0] = 16'hFF99	;
     501: sin_wave[15:0] = 16'hFECB	;
     502: sin_wave[15:0] = 16'hFDFD	;
     503: sin_wave[15:0] = 16'hFD2F	;
     504: sin_wave[15:0] = 16'hFC61	;
     505: sin_wave[15:0] = 16'hFB93	;
     506: sin_wave[15:0] = 16'hFAC5	;
     507: sin_wave[15:0] = 16'hF9F7	;
     508: sin_wave[15:0] = 16'hF929	;
     509: sin_wave[15:0] = 16'hF85B	;
     510: sin_wave[15:0] = 16'hF78E	;
     511: sin_wave[15:0] = 16'hF6C0	;
     512: sin_wave[15:0] = 16'hF5F3	;
     513: sin_wave[15:0] = 16'hF525	;
     514: sin_wave[15:0] = 16'hF458	;
     515: sin_wave[15:0] = 16'hF38B	;
     516: sin_wave[15:0] = 16'hF2BE	;
     517: sin_wave[15:0] = 16'hF1F1	;
     518: sin_wave[15:0] = 16'hF124	;
     519: sin_wave[15:0] = 16'hF057	;
     520: sin_wave[15:0] = 16'hEF8B	;
     521: sin_wave[15:0] = 16'hEEBF	;
     522: sin_wave[15:0] = 16'hEDF2	;
     523: sin_wave[15:0] = 16'hED27	;
     524: sin_wave[15:0] = 16'hEC5B	;
     525: sin_wave[15:0] = 16'hEB8F	;
     526: sin_wave[15:0] = 16'hEAC4	;
     527: sin_wave[15:0] = 16'hE9F9	;
     528: sin_wave[15:0] = 16'hE92E	;
     529: sin_wave[15:0] = 16'hE863	;
     530: sin_wave[15:0] = 16'hE799	;
     531: sin_wave[15:0] = 16'hE6CF	;
     532: sin_wave[15:0] = 16'hE605	;
     533: sin_wave[15:0] = 16'hE53B	;
     534: sin_wave[15:0] = 16'hE472	;
     535: sin_wave[15:0] = 16'hE3A9	;
     536: sin_wave[15:0] = 16'hE2E0	;
     537: sin_wave[15:0] = 16'hE217	;
     538: sin_wave[15:0] = 16'hE14F	;
     539: sin_wave[15:0] = 16'hE087	;
     540: sin_wave[15:0] = 16'hDFBF	;
     541: sin_wave[15:0] = 16'hDEF8	;
     542: sin_wave[15:0] = 16'hDE31	;
     543: sin_wave[15:0] = 16'hDD6B	;
     544: sin_wave[15:0] = 16'hDCA4	;
     545: sin_wave[15:0] = 16'hDBDE	;
     546: sin_wave[15:0] = 16'hDB19	;
     547: sin_wave[15:0] = 16'hDA54	;
     548: sin_wave[15:0] = 16'hD98F	;
     549: sin_wave[15:0] = 16'hD8CB	;
     550: sin_wave[15:0] = 16'hD807	;
     551: sin_wave[15:0] = 16'hD743	;
     552: sin_wave[15:0] = 16'hD680	;
     553: sin_wave[15:0] = 16'hD5BD	;
     554: sin_wave[15:0] = 16'hD4FB	;
     555: sin_wave[15:0] = 16'hD439	;
     556: sin_wave[15:0] = 16'hD378	;
     557: sin_wave[15:0] = 16'hD2B7	;
     558: sin_wave[15:0] = 16'hD1F6	;
     559: sin_wave[15:0] = 16'hD136	;
     560: sin_wave[15:0] = 16'hD076	;
     561: sin_wave[15:0] = 16'hCFB7	;
     562: sin_wave[15:0] = 16'hCEF9	;
     563: sin_wave[15:0] = 16'hCE3B	;
     564: sin_wave[15:0] = 16'hCD7D	;
     565: sin_wave[15:0] = 16'hCCC0	;
     566: sin_wave[15:0] = 16'hCC03	;
     567: sin_wave[15:0] = 16'hCB47	;
     568: sin_wave[15:0] = 16'hCA8C	;
     569: sin_wave[15:0] = 16'hC9D1	;
     570: sin_wave[15:0] = 16'hC916	;
     571: sin_wave[15:0] = 16'hC85C	;
     572: sin_wave[15:0] = 16'hC7A3	;
     573: sin_wave[15:0] = 16'hC6EA	;
     574: sin_wave[15:0] = 16'hC632	;
     575: sin_wave[15:0] = 16'hC57B	;
     576: sin_wave[15:0] = 16'hC4C4	;
     577: sin_wave[15:0] = 16'hC40D	;
     578: sin_wave[15:0] = 16'hC357	;
     579: sin_wave[15:0] = 16'hC2A2	;
     580: sin_wave[15:0] = 16'hC1EE	;
     581: sin_wave[15:0] = 16'hC13A	;
     582: sin_wave[15:0] = 16'hC087	;
     583: sin_wave[15:0] = 16'hBFD4	;
     584: sin_wave[15:0] = 16'hBF22	;
     585: sin_wave[15:0] = 16'hBE71	;
     586: sin_wave[15:0] = 16'hBDC0	;
     587: sin_wave[15:0] = 16'hBD10	;
     588: sin_wave[15:0] = 16'hBC61	;
     589: sin_wave[15:0] = 16'hBBB2	;
     590: sin_wave[15:0] = 16'hBB04	;
     591: sin_wave[15:0] = 16'hBA57	;
     592: sin_wave[15:0] = 16'hB9AA	;
     593: sin_wave[15:0] = 16'hB8FE	;
     594: sin_wave[15:0] = 16'hB853	;
     595: sin_wave[15:0] = 16'hB7A9	;
     596: sin_wave[15:0] = 16'hB6FF	;
     597: sin_wave[15:0] = 16'hB656	;
     598: sin_wave[15:0] = 16'hB5AE	;
     599: sin_wave[15:0] = 16'hB507	;
     600: sin_wave[15:0] = 16'hB460	;
     601: sin_wave[15:0] = 16'hB3BA	;
     602: sin_wave[15:0] = 16'hB315	;
     603: sin_wave[15:0] = 16'hB271	;
     604: sin_wave[15:0] = 16'hB1CD	;
     605: sin_wave[15:0] = 16'hB12B	;
     606: sin_wave[15:0] = 16'hB089	;
     607: sin_wave[15:0] = 16'hAFE7	;
     608: sin_wave[15:0] = 16'hAF47	;
     609: sin_wave[15:0] = 16'hAEA8	;
     610: sin_wave[15:0] = 16'hAE09	;
     611: sin_wave[15:0] = 16'hAD6B	;
     612: sin_wave[15:0] = 16'hACCE	;
     613: sin_wave[15:0] = 16'hAC32	;
     614: sin_wave[15:0] = 16'hAB96	;
     615: sin_wave[15:0] = 16'hAAFC	;
     616: sin_wave[15:0] = 16'hAA62	;
     617: sin_wave[15:0] = 16'hA9C9	;
     618: sin_wave[15:0] = 16'hA932	;
     619: sin_wave[15:0] = 16'hA89B	;
     620: sin_wave[15:0] = 16'hA804	;
     621: sin_wave[15:0] = 16'hA76F	;
     622: sin_wave[15:0] = 16'hA6DB	;
     623: sin_wave[15:0] = 16'hA647	;
     624: sin_wave[15:0] = 16'hA5B5	;
     625: sin_wave[15:0] = 16'hA523	;
     626: sin_wave[15:0] = 16'hA493	;
     627: sin_wave[15:0] = 16'hA403	;
     628: sin_wave[15:0] = 16'hA374	;
     629: sin_wave[15:0] = 16'hA2E6	;
     630: sin_wave[15:0] = 16'hA259	;
     631: sin_wave[15:0] = 16'hA1CD	;
     632: sin_wave[15:0] = 16'hA142	;
     633: sin_wave[15:0] = 16'hA0B8	;
     634: sin_wave[15:0] = 16'hA02F	;
     635: sin_wave[15:0] = 16'h9FA7	;
     636: sin_wave[15:0] = 16'h9F20	;
     637: sin_wave[15:0] = 16'h9E99	;
     638: sin_wave[15:0] = 16'h9E14	;
     639: sin_wave[15:0] = 16'h9D90	;
     640: sin_wave[15:0] = 16'h9D0D	;
     641: sin_wave[15:0] = 16'h9C8B	;
     642: sin_wave[15:0] = 16'h9C09	;
     643: sin_wave[15:0] = 16'h9B89	;
     644: sin_wave[15:0] = 16'h9B0A	;
     645: sin_wave[15:0] = 16'h9A8C	;
     646: sin_wave[15:0] = 16'h9A0F	;
     647: sin_wave[15:0] = 16'h9992	;
     648: sin_wave[15:0] = 16'h9917	;
     649: sin_wave[15:0] = 16'h989D	;
     650: sin_wave[15:0] = 16'h9824	;
     651: sin_wave[15:0] = 16'h97AC	;
     652: sin_wave[15:0] = 16'h9736	;
     653: sin_wave[15:0] = 16'h96C0	;
     654: sin_wave[15:0] = 16'h964B	;
     655: sin_wave[15:0] = 16'h95D7	;
     656: sin_wave[15:0] = 16'h9565	;
     657: sin_wave[15:0] = 16'h94F3	;
     658: sin_wave[15:0] = 16'h9483	;
     659: sin_wave[15:0] = 16'h9414	;
     660: sin_wave[15:0] = 16'h93A5	;
     661: sin_wave[15:0] = 16'h9338	;
     662: sin_wave[15:0] = 16'h92CC	;
     663: sin_wave[15:0] = 16'h9261	;
     664: sin_wave[15:0] = 16'h91F7	;
     665: sin_wave[15:0] = 16'h918F	;
     666: sin_wave[15:0] = 16'h9127	;
     667: sin_wave[15:0] = 16'h90C0	;
     668: sin_wave[15:0] = 16'h905B	;
     669: sin_wave[15:0] = 16'h8FF7	;
     670: sin_wave[15:0] = 16'h8F94	;
     671: sin_wave[15:0] = 16'h8F32	;
     672: sin_wave[15:0] = 16'h8ED1	;
     673: sin_wave[15:0] = 16'h8E71	;
     674: sin_wave[15:0] = 16'h8E13	;
     675: sin_wave[15:0] = 16'h8DB5	;
     676: sin_wave[15:0] = 16'h8D59	;
     677: sin_wave[15:0] = 16'h8CFE	;
     678: sin_wave[15:0] = 16'h8CA4	;
     679: sin_wave[15:0] = 16'h8C4C	;
     680: sin_wave[15:0] = 16'h8BF4	;
     681: sin_wave[15:0] = 16'h8B9E	;
     682: sin_wave[15:0] = 16'h8B49	;
     683: sin_wave[15:0] = 16'h8AF5	;
     684: sin_wave[15:0] = 16'h8AA2	;
     685: sin_wave[15:0] = 16'h8A50	;
     686: sin_wave[15:0] = 16'h8A00	;
     687: sin_wave[15:0] = 16'h89B0	;
     688: sin_wave[15:0] = 16'h8962	;
     689: sin_wave[15:0] = 16'h8916	;
     690: sin_wave[15:0] = 16'h88CA	;
     691: sin_wave[15:0] = 16'h8880	;
     692: sin_wave[15:0] = 16'h8836	;
     693: sin_wave[15:0] = 16'h87EE	;
     694: sin_wave[15:0] = 16'h87A8	;
     695: sin_wave[15:0] = 16'h8762	;
     696: sin_wave[15:0] = 16'h871E	;
     697: sin_wave[15:0] = 16'h86DA	;
     698: sin_wave[15:0] = 16'h8699	;
     699: sin_wave[15:0] = 16'h8658	;
     700: sin_wave[15:0] = 16'h8618	;
     701: sin_wave[15:0] = 16'h85DA	;
     702: sin_wave[15:0] = 16'h859D	;
     703: sin_wave[15:0] = 16'h8562	;
     704: sin_wave[15:0] = 16'h8527	;
     705: sin_wave[15:0] = 16'h84EE	;
     706: sin_wave[15:0] = 16'h84B6	;
     707: sin_wave[15:0] = 16'h847F	;
     708: sin_wave[15:0] = 16'h844A	;
     709: sin_wave[15:0] = 16'h8415	;
     710: sin_wave[15:0] = 16'h83E2	;
     711: sin_wave[15:0] = 16'h83B1	;
     712: sin_wave[15:0] = 16'h8380	;
     713: sin_wave[15:0] = 16'h8351	;
     714: sin_wave[15:0] = 16'h8323	;
     715: sin_wave[15:0] = 16'h82F6	;
     716: sin_wave[15:0] = 16'h82CB	;
     717: sin_wave[15:0] = 16'h82A1	;
     718: sin_wave[15:0] = 16'h8278	;
     719: sin_wave[15:0] = 16'h8250	;
     720: sin_wave[15:0] = 16'h822A	;
     721: sin_wave[15:0] = 16'h8205	;
     722: sin_wave[15:0] = 16'h81E1	;
     723: sin_wave[15:0] = 16'h81BF	;
     724: sin_wave[15:0] = 16'h819D	;
     725: sin_wave[15:0] = 16'h817D	;
     726: sin_wave[15:0] = 16'h815F	;
     727: sin_wave[15:0] = 16'h8141	;
     728: sin_wave[15:0] = 16'h8125	;
     729: sin_wave[15:0] = 16'h810A	;
     730: sin_wave[15:0] = 16'h80F1	;
     731: sin_wave[15:0] = 16'h80D9	;
     732: sin_wave[15:0] = 16'h80C2	;
     733: sin_wave[15:0] = 16'h80AC	;
     734: sin_wave[15:0] = 16'h8098	;
     735: sin_wave[15:0] = 16'h8085	;
     736: sin_wave[15:0] = 16'h8073	;
     737: sin_wave[15:0] = 16'h8062	;
     738: sin_wave[15:0] = 16'h8053	;
     739: sin_wave[15:0] = 16'h8045	;
     740: sin_wave[15:0] = 16'h8038	;
     741: sin_wave[15:0] = 16'h802D	;
     742: sin_wave[15:0] = 16'h8023	;
     743: sin_wave[15:0] = 16'h801A	;
     744: sin_wave[15:0] = 16'h8013	;
     745: sin_wave[15:0] = 16'h800D	;
     746: sin_wave[15:0] = 16'h8008	;
     747: sin_wave[15:0] = 16'h8004	;
     748: sin_wave[15:0] = 16'h8002	;
     749: sin_wave[15:0] = 16'h8001	;
     750: sin_wave[15:0] = 16'h8001	;
     751: sin_wave[15:0] = 16'h8003	;
     752: sin_wave[15:0] = 16'h8006	;
     753: sin_wave[15:0] = 16'h800A	;
     754: sin_wave[15:0] = 16'h8010	;
     755: sin_wave[15:0] = 16'h8016	;
     756: sin_wave[15:0] = 16'h801F	;
     757: sin_wave[15:0] = 16'h8028	;
     758: sin_wave[15:0] = 16'h8033	;
     759: sin_wave[15:0] = 16'h803F	;
     760: sin_wave[15:0] = 16'h804C	;
     761: sin_wave[15:0] = 16'h805A	;
     762: sin_wave[15:0] = 16'h806A	;
     763: sin_wave[15:0] = 16'h807B	;
     764: sin_wave[15:0] = 16'h808E	;
     765: sin_wave[15:0] = 16'h80A2	;
     766: sin_wave[15:0] = 16'h80B7	;
     767: sin_wave[15:0] = 16'h80CD	;
     768: sin_wave[15:0] = 16'h80E5	;
     769: sin_wave[15:0] = 16'h80FD	;
     770: sin_wave[15:0] = 16'h8118	;
     771: sin_wave[15:0] = 16'h8133	;
     772: sin_wave[15:0] = 16'h8150	;
     773: sin_wave[15:0] = 16'h816E	;
     774: sin_wave[15:0] = 16'h818D	;
     775: sin_wave[15:0] = 16'h81AE	;
     776: sin_wave[15:0] = 16'h81D0	;
     777: sin_wave[15:0] = 16'h81F3	;
     778: sin_wave[15:0] = 16'h8217	;
     779: sin_wave[15:0] = 16'h823D	;
     780: sin_wave[15:0] = 16'h8264	;
     781: sin_wave[15:0] = 16'h828C	;
     782: sin_wave[15:0] = 16'h82B6	;
     783: sin_wave[15:0] = 16'h82E0	;
     784: sin_wave[15:0] = 16'h830C	;
     785: sin_wave[15:0] = 16'h833A	;
     786: sin_wave[15:0] = 16'h8368	;
     787: sin_wave[15:0] = 16'h8398	;
     788: sin_wave[15:0] = 16'h83C9	;
     789: sin_wave[15:0] = 16'h83FC	;
     790: sin_wave[15:0] = 16'h842F	;
     791: sin_wave[15:0] = 16'h8464	;
     792: sin_wave[15:0] = 16'h849A	;
     793: sin_wave[15:0] = 16'h84D2	;
     794: sin_wave[15:0] = 16'h850A	;
     795: sin_wave[15:0] = 16'h8544	;
     796: sin_wave[15:0] = 16'h857F	;
     797: sin_wave[15:0] = 16'h85BC	;
     798: sin_wave[15:0] = 16'h85F9	;
     799: sin_wave[15:0] = 16'h8638	;
     800: sin_wave[15:0] = 16'h8678	;
     801: sin_wave[15:0] = 16'h86B9	;
     802: sin_wave[15:0] = 16'h86FC	;
     803: sin_wave[15:0] = 16'h8740	;
     804: sin_wave[15:0] = 16'h8785	;
     805: sin_wave[15:0] = 16'h87CB	;
     806: sin_wave[15:0] = 16'h8812	;
     807: sin_wave[15:0] = 16'h885B	;
     808: sin_wave[15:0] = 16'h88A5	;
     809: sin_wave[15:0] = 16'h88F0	;
     810: sin_wave[15:0] = 16'h893C	;
     811: sin_wave[15:0] = 16'h8989	;
     812: sin_wave[15:0] = 16'h89D8	;
     813: sin_wave[15:0] = 16'h8A28	;
     814: sin_wave[15:0] = 16'h8A79	;
     815: sin_wave[15:0] = 16'h8ACB	;
     816: sin_wave[15:0] = 16'h8B1E	;
     817: sin_wave[15:0] = 16'h8B73	;
     818: sin_wave[15:0] = 16'h8BC9	;
     819: sin_wave[15:0] = 16'h8C20	;
     820: sin_wave[15:0] = 16'h8C78	;
     821: sin_wave[15:0] = 16'h8CD1	;
     822: sin_wave[15:0] = 16'h8D2C	;
     823: sin_wave[15:0] = 16'h8D87	;
     824: sin_wave[15:0] = 16'h8DE4	;
     825: sin_wave[15:0] = 16'h8E42	;
     826: sin_wave[15:0] = 16'h8EA1	;
     827: sin_wave[15:0] = 16'h8F01	;
     828: sin_wave[15:0] = 16'h8F63	;
     829: sin_wave[15:0] = 16'h8FC5	;
     830: sin_wave[15:0] = 16'h9029	;
     831: sin_wave[15:0] = 16'h908E	;
     832: sin_wave[15:0] = 16'h90F4	;
     833: sin_wave[15:0] = 16'h915B	;
     834: sin_wave[15:0] = 16'h91C3	;
     835: sin_wave[15:0] = 16'h922C	;
     836: sin_wave[15:0] = 16'h9296	;
     837: sin_wave[15:0] = 16'h9302	;
     838: sin_wave[15:0] = 16'h936F	;
     839: sin_wave[15:0] = 16'h93DC	;
     840: sin_wave[15:0] = 16'h944B	;
     841: sin_wave[15:0] = 16'h94BB	;
     842: sin_wave[15:0] = 16'h952C	;
     843: sin_wave[15:0] = 16'h959E	;
     844: sin_wave[15:0] = 16'h9611	;
     845: sin_wave[15:0] = 16'h9685	;
     846: sin_wave[15:0] = 16'h96FB	;
     847: sin_wave[15:0] = 16'h9771	;
     848: sin_wave[15:0] = 16'h97E8	;
     849: sin_wave[15:0] = 16'h9861	;
     850: sin_wave[15:0] = 16'h98DA	;
     851: sin_wave[15:0] = 16'h9955	;
     852: sin_wave[15:0] = 16'h99D0	;
     853: sin_wave[15:0] = 16'h9A4D	;
     854: sin_wave[15:0] = 16'h9ACB	;
     855: sin_wave[15:0] = 16'h9B49	;
     856: sin_wave[15:0] = 16'h9BC9	;
     857: sin_wave[15:0] = 16'h9C4A	;
     858: sin_wave[15:0] = 16'h9CCB	;
     859: sin_wave[15:0] = 16'h9D4E	;
     860: sin_wave[15:0] = 16'h9DD2	;
     861: sin_wave[15:0] = 16'h9E57	;
     862: sin_wave[15:0] = 16'h9EDC	;
     863: sin_wave[15:0] = 16'h9F63	;
     864: sin_wave[15:0] = 16'h9FEB	;
     865: sin_wave[15:0] = 16'hA073	;
     866: sin_wave[15:0] = 16'hA0FD	;
     867: sin_wave[15:0] = 16'hA188	;
     868: sin_wave[15:0] = 16'hA213	;
     869: sin_wave[15:0] = 16'hA2A0	;
     870: sin_wave[15:0] = 16'hA32D	;
     871: sin_wave[15:0] = 16'hA3BB	;
     872: sin_wave[15:0] = 16'hA44B	;
     873: sin_wave[15:0] = 16'hA4DB	;
     874: sin_wave[15:0] = 16'hA56C	;
     875: sin_wave[15:0] = 16'hA5FE	;
     876: sin_wave[15:0] = 16'hA691	;
     877: sin_wave[15:0] = 16'hA725	;
     878: sin_wave[15:0] = 16'hA7BA	;
     879: sin_wave[15:0] = 16'hA84F	;
     880: sin_wave[15:0] = 16'hA8E6	;
     881: sin_wave[15:0] = 16'hA97D	;
     882: sin_wave[15:0] = 16'hAA16	;
     883: sin_wave[15:0] = 16'hAAAF	;
     884: sin_wave[15:0] = 16'hAB49	;
     885: sin_wave[15:0] = 16'hABE4	;
     886: sin_wave[15:0] = 16'hAC80	;
     887: sin_wave[15:0] = 16'hAD1C	;
     888: sin_wave[15:0] = 16'hADBA	;
     889: sin_wave[15:0] = 16'hAE58	;
     890: sin_wave[15:0] = 16'hAEF7	;
     891: sin_wave[15:0] = 16'hAF97	;
     892: sin_wave[15:0] = 16'hB038	;
     893: sin_wave[15:0] = 16'hB0D9	;
     894: sin_wave[15:0] = 16'hB17C	;
     895: sin_wave[15:0] = 16'hB21F	;
     896: sin_wave[15:0] = 16'hB2C3	;
     897: sin_wave[15:0] = 16'hB368	;
     898: sin_wave[15:0] = 16'hB40D	;
     899: sin_wave[15:0] = 16'hB4B3	;
     900: sin_wave[15:0] = 16'hB55A	;
     901: sin_wave[15:0] = 16'hB602	;
     902: sin_wave[15:0] = 16'hB6AB	;
     903: sin_wave[15:0] = 16'hB754	;
     904: sin_wave[15:0] = 16'hB7FE	;
     905: sin_wave[15:0] = 16'hB8A9	;
     906: sin_wave[15:0] = 16'hB954	;
     907: sin_wave[15:0] = 16'hBA00	;
     908: sin_wave[15:0] = 16'hBAAD	;
     909: sin_wave[15:0] = 16'hBB5B	;
     910: sin_wave[15:0] = 16'hBC09	;
     911: sin_wave[15:0] = 16'hBCB8	;
     912: sin_wave[15:0] = 16'hBD68	;
     913: sin_wave[15:0] = 16'hBE18	;
     914: sin_wave[15:0] = 16'hBEC9	;
     915: sin_wave[15:0] = 16'hBF7B	;
     916: sin_wave[15:0] = 16'hC02D	;
     917: sin_wave[15:0] = 16'hC0E0	;
     918: sin_wave[15:0] = 16'hC194	;
     919: sin_wave[15:0] = 16'hC248	;
     920: sin_wave[15:0] = 16'hC2FD	;
     921: sin_wave[15:0] = 16'hC3B2	;
     922: sin_wave[15:0] = 16'hC468	;
     923: sin_wave[15:0] = 16'hC51F	;
     924: sin_wave[15:0] = 16'hC5D6	;
     925: sin_wave[15:0] = 16'hC68E	;
     926: sin_wave[15:0] = 16'hC747	;
     927: sin_wave[15:0] = 16'hC800	;
     928: sin_wave[15:0] = 16'hC8B9	;
     929: sin_wave[15:0] = 16'hC973	;
     930: sin_wave[15:0] = 16'hCA2E	;
     931: sin_wave[15:0] = 16'hCAE9	;
     932: sin_wave[15:0] = 16'hCBA5	;
     933: sin_wave[15:0] = 16'hCC62	;
     934: sin_wave[15:0] = 16'hCD1E	;
     935: sin_wave[15:0] = 16'hCDDC	;
     936: sin_wave[15:0] = 16'hCE9A	;
     937: sin_wave[15:0] = 16'hCF58	;
     938: sin_wave[15:0] = 16'hD017	;
     939: sin_wave[15:0] = 16'hD0D6	;
     940: sin_wave[15:0] = 16'hD196	;
     941: sin_wave[15:0] = 16'hD256	;
     942: sin_wave[15:0] = 16'hD317	;
     943: sin_wave[15:0] = 16'hD3D8	;
     944: sin_wave[15:0] = 16'hD49A	;
     945: sin_wave[15:0] = 16'hD55C	;
     946: sin_wave[15:0] = 16'hD61F	;
     947: sin_wave[15:0] = 16'hD6E1	;
     948: sin_wave[15:0] = 16'hD7A5	;
     949: sin_wave[15:0] = 16'hD869	;
     950: sin_wave[15:0] = 16'hD92D	;
     951: sin_wave[15:0] = 16'hD9F1	;
     952: sin_wave[15:0] = 16'hDAB6	;
     953: sin_wave[15:0] = 16'hDB7C	;
     954: sin_wave[15:0] = 16'hDC41	;
     955: sin_wave[15:0] = 16'hDD07	;
     956: sin_wave[15:0] = 16'hDDCE	;
     957: sin_wave[15:0] = 16'hDE95	;
     958: sin_wave[15:0] = 16'hDF5C	;
     959: sin_wave[15:0] = 16'hE023	;
     960: sin_wave[15:0] = 16'hE0EB	;
     961: sin_wave[15:0] = 16'hE1B3	;
     962: sin_wave[15:0] = 16'hE27B	;
     963: sin_wave[15:0] = 16'hE344	;
     964: sin_wave[15:0] = 16'hE40D	;
     965: sin_wave[15:0] = 16'hE4D6	;
     966: sin_wave[15:0] = 16'hE5A0	;
     967: sin_wave[15:0] = 16'hE66A	;
     968: sin_wave[15:0] = 16'hE734	;
     969: sin_wave[15:0] = 16'hE7FE	;
     970: sin_wave[15:0] = 16'hE8C9	;
     971: sin_wave[15:0] = 16'hE993	;
     972: sin_wave[15:0] = 16'hEA5E	;
     973: sin_wave[15:0] = 16'hEB2A	;
     974: sin_wave[15:0] = 16'hEBF5	;
     975: sin_wave[15:0] = 16'hECC1	;
     976: sin_wave[15:0] = 16'hED8D	;
     977: sin_wave[15:0] = 16'hEE59	;
     978: sin_wave[15:0] = 16'hEF25	;
     979: sin_wave[15:0] = 16'hEFF1	;
     980: sin_wave[15:0] = 16'hF0BE	;
     981: sin_wave[15:0] = 16'hF18A	;
     982: sin_wave[15:0] = 16'hF257	;
     983: sin_wave[15:0] = 16'hF324	;
     984: sin_wave[15:0] = 16'hF3F1	;
     985: sin_wave[15:0] = 16'hF4BF	;
     986: sin_wave[15:0] = 16'hF58C	;
     987: sin_wave[15:0] = 16'hF659	;
     988: sin_wave[15:0] = 16'hF727	;
     989: sin_wave[15:0] = 16'hF7F4	;
     990: sin_wave[15:0] = 16'hF8C2	;
     991: sin_wave[15:0] = 16'hF990	;
     992: sin_wave[15:0] = 16'hFA5E	;
     993: sin_wave[15:0] = 16'hFB2C	;
     994: sin_wave[15:0] = 16'hFBFA	;
     995: sin_wave[15:0] = 16'hFCC8	;
     996: sin_wave[15:0] = 16'hFD96	;
     997: sin_wave[15:0] = 16'hFE64	;
     998: sin_wave[15:0] = 16'hFF32	;
     999: sin_wave[15:0] = 16'h0000	;
     endcase
end
//    
endmodule
